// $Id$
// ncgen -b -o ${DATA}/aca/idx_rfr_roush_montmorillonite.nc ${HOME}/idx_rfr/idx_rfr_roush_montmorillonite.cdl

netcdf idx_rfr_roush_montmorillonite {

dimensions:
	bnd = 401 ;

variables:

// global attributes:
	:RCS_Header = "$Id$" ;
	:history = "" ;
	:description = "Montmorillonite refractive indices" ;
	:source="
T. Roush (NASA Ames), Pollack, and Orenberg Icarus 94, 1991
Ultimate source is T. Roush (NASA Ames)
Brian Hansell (UCLA) converted data from T. Roush into netCDF format 01 October, 2005.
Charlie Zender (zender at uci dot edu) standardized 20060129.
	";

	float bnd(bnd) ;
		bnd:units = "microns" ;
		bnd:longname = "band center wavelength" ;
		bnd:C_format = "%.5g" ;

	float idx_rfr_montmorillonite_rl(bnd) ;
		idx_rfr_montmorillonite_rl:units = "" ;
		idx_rfr_montmorillonite_rl:longname = "Montmorillonite refractive index, real" ;
		idx_rfr_montmorillonite_rl:C_format = "%.4g" ;

	float idx_rfr_montmorillonite_img(bnd) ;
		idx_rfr_montmorillonite_img:units = "" ;
		idx_rfr_montmorillonite_img:longname = "Montmorillonite refractive index, imaginary" ;
		idx_rfr_montmorillonite_img:C_format = "%.3g" ;

data:

 bnd = 5, 5.01, 5.02, 5.03, 5.04, 5.05, 5.061, 5.071, 5.081, 5.092, 5.102, 
    5.113, 5.123, 5.134, 5.144, 5.155, 5.165, 5.176, 5.187, 5.198, 5.208, 
    5.219, 5.23, 5.241, 5.252, 5.263, 5.274, 5.285, 5.297, 5.308, 5.319, 
    5.331, 5.342, 5.353, 5.365, 5.376, 5.388, 5.4, 5.411, 5.423, 5.435, 
    5.447, 5.458, 5.47, 5.483, 5.495, 5.507, 5.519, 5.531, 5.543, 5.556, 
    5.568, 5.58, 5.593, 5.605, 5.618, 5.631, 5.643, 5.656, 5.669, 5.682, 
    5.695, 5.708, 5.721, 5.734, 5.747, 5.76, 5.774, 5.787, 5.8, 5.814, 5.827, 
    5.841, 5.855, 5.869, 5.882, 5.896, 5.91, 5.924, 5.938, 5.952, 5.967, 
    5.981, 5.995, 6.01, 6.024, 6.039, 6.053, 6.068, 6.083, 6.098, 6.113, 
    6.128, 6.142, 6.158, 6.173, 6.188, 6.203, 6.219, 6.234, 6.25, 6.266, 
    6.281, 6.297, 6.313, 6.329, 6.345, 6.361, 6.378, 6.394, 6.41, 6.427, 
    6.443, 6.46, 6.477, 6.494, 6.51, 6.527, 6.544, 6.562, 6.579, 6.596, 
    6.614, 6.631, 6.649, 6.667, 6.685, 6.702, 6.72, 6.739, 6.757, 6.775, 
    6.793, 6.812, 6.831, 6.849, 6.868, 6.887, 6.906, 6.925, 6.944, 6.964, 
    6.983, 7.003, 7.023, 7.042, 7.062, 7.082, 7.102, 7.122, 7.143, 7.163, 
    7.184, 7.205, 7.225, 7.246, 7.267, 7.289, 7.31, 7.331, 7.353, 7.375, 
    7.396, 7.418, 7.44, 7.463, 7.485, 7.508, 7.53, 7.553, 7.576, 7.599, 
    7.622, 7.645, 7.669, 7.692, 7.716, 7.74, 7.764, 7.788, 7.813, 7.837, 
    7.862, 7.886, 7.911, 7.937, 7.962, 7.987, 8.013, 8.039, 8.064, 8.091, 
    8.117, 8.143, 8.17, 8.197, 8.224, 8.251, 8.278, 8.306, 8.333, 8.361, 
    8.389, 8.417, 8.446, 8.475, 8.503, 8.532, 8.562, 8.591, 8.621, 8.651, 
    8.681, 8.711, 8.741, 8.772, 8.803, 8.834, 8.865, 8.897, 8.929, 8.961, 
    8.993, 9.025, 9.058, 9.091, 9.124, 9.158, 9.191, 9.225, 9.259, 9.294, 
    9.328, 9.363, 9.399, 9.434, 9.47, 9.506, 9.542, 9.578, 9.615, 9.653, 
    9.69, 9.728, 9.766, 9.804, 9.842, 9.881, 9.921, 9.96, 10, 10.04, 10.081, 
    10.121, 10.163, 10.204, 10.246, 10.288, 10.331, 10.373, 10.417, 10.46, 
    10.504, 10.549, 10.593, 10.638, 10.684, 10.73, 10.776, 10.823, 10.87, 
    10.917, 10.965, 11.013, 11.062, 11.111, 11.161, 11.211, 11.261, 11.312, 
    11.364, 11.416, 11.468, 11.521, 11.574, 11.628, 11.682, 11.737, 11.792, 
    11.848, 11.905, 11.962, 12.019, 12.077, 12.136, 12.195, 12.255, 12.315, 
    12.376, 12.438, 12.5, 12.563, 12.626, 12.69, 12.755, 12.821, 12.887, 
    12.953, 13.021, 13.089, 13.158, 13.228, 13.298, 13.369, 13.441, 13.514, 
    13.587, 13.661, 13.736, 13.812, 13.889, 13.966, 14.045, 14.124, 14.205, 
    14.286, 14.368, 14.451, 14.535, 14.62, 14.706, 14.793, 14.881, 14.97, 
    15.06, 15.152, 15.244, 15.337, 15.432, 15.528, 15.625, 15.723, 15.823, 
    15.924, 16.026, 16.129, 16.234, 16.34, 16.447, 16.556, 16.667, 16.779, 
    16.892, 17.007, 17.123, 17.241, 17.361, 17.483, 17.606, 17.731, 17.857, 
    17.986, 18.116, 18.248, 18.382, 18.519, 18.657, 18.797, 18.939, 19.084, 
    19.231, 19.38, 19.531, 19.685, 19.841, 20, 20.161, 20.325, 20.492, 
    20.661, 20.833, 21.008, 21.186, 21.368, 21.552, 21.739, 21.93, 22.124, 
    22.321, 22.523, 22.727, 22.936, 23.148, 23.364, 23.585, 23.81, 24.038, 
    24.272, 24.51, 24.752, 25 ;

 idx_rfr_montmorillonite_rl = 1.336, 1.335, 1.335, 1.335, 1.334, 1.334, 
    1.333, 1.333, 1.333, 1.332, 1.332, 1.332, 1.331, 1.331, 1.33, 1.33, 
    1.329, 1.329, 1.329, 1.328, 1.328, 1.327, 1.327, 1.326, 1.326, 1.325, 
    1.325, 1.324, 1.324, 1.324, 1.323, 1.322, 1.322, 1.321, 1.321, 1.32, 
    1.32, 1.319, 1.319, 1.318, 1.318, 1.317, 1.317, 1.316, 1.316, 1.315, 
    1.314, 1.314, 1.313, 1.313, 1.312, 1.311, 1.311, 1.31, 1.309, 1.309, 
    1.308, 1.308, 1.307, 1.306, 1.305, 1.305, 1.304, 1.303, 1.302, 1.302, 
    1.301, 1.3, 1.299, 1.298, 1.298, 1.297, 1.296, 1.295, 1.294, 1.293, 
    1.292, 1.291, 1.29, 1.289, 1.288, 1.287, 1.285, 1.284, 1.282, 1.281, 
    1.279, 1.276, 1.274, 1.271, 1.269, 1.272, 1.284, 1.294, 1.294, 1.291, 
    1.288, 1.286, 1.283, 1.281, 1.28, 1.278, 1.276, 1.275, 1.273, 1.271, 
    1.27, 1.269, 1.267, 1.266, 1.264, 1.263, 1.261, 1.26, 1.258, 1.257, 
    1.256, 1.254, 1.253, 1.251, 1.25, 1.248, 1.246, 1.245, 1.243, 1.241, 
    1.24, 1.238, 1.236, 1.234, 1.232, 1.231, 1.229, 1.227, 1.225, 1.223, 
    1.221, 1.219, 1.217, 1.214, 1.212, 1.21, 1.208, 1.205, 1.203, 1.201, 
    1.198, 1.195, 1.193, 1.19, 1.187, 1.185, 1.182, 1.179, 1.176, 1.173, 
    1.169, 1.166, 1.163, 1.159, 1.156, 1.152, 1.148, 1.145, 1.141, 1.137, 
    1.132, 1.128, 1.124, 1.119, 1.114, 1.109, 1.104, 1.099, 1.094, 1.088, 
    1.082, 1.076, 1.07, 1.063, 1.056, 1.049, 1.042, 1.034, 1.026, 1.018, 
    1.009, 1, 0.99, 0.98, 0.969, 0.957, 0.945, 0.933, 0.919, 0.905, 0.89, 
    0.874, 0.856, 0.838, 0.818, 0.797, 0.774, 0.75, 0.725, 0.699, 0.672, 
    0.645, 0.621, 0.6, 0.585, 0.577, 0.575, 0.579, 0.587, 0.601, 0.625, 
    0.663, 0.716, 0.777, 0.826, 0.844, 0.824, 0.779, 0.724, 0.671, 0.63, 
    0.605, 0.598, 0.609, 0.637, 0.684, 0.754, 0.851, 0.982, 1.153, 1.365, 
    1.601, 1.823, 1.986, 2.078, 2.126, 2.177, 2.259, 2.365, 2.458, 2.504, 
    2.501, 2.464, 2.409, 2.349, 2.289, 2.232, 2.179, 2.129, 2.084, 2.042, 
    2.003, 1.966, 1.932, 1.899, 1.868, 1.838, 1.809, 1.78, 1.752, 1.726, 
    1.706, 1.698, 1.713, 1.748, 1.777, 1.782, 1.769, 1.749, 1.727, 1.707, 
    1.692, 1.688, 1.695, 1.704, 1.705, 1.697, 1.682, 1.665, 1.648, 1.637, 
    1.642, 1.648, 1.639, 1.624, 1.61, 1.596, 1.583, 1.57, 1.558, 1.546, 
    1.533, 1.521, 1.51, 1.503, 1.505, 1.517, 1.527, 1.526, 1.518, 1.507, 
    1.495, 1.484, 1.474, 1.463, 1.453, 1.443, 1.433, 1.423, 1.412, 1.402, 
    1.392, 1.381, 1.37, 1.359, 1.347, 1.335, 1.323, 1.313, 1.308, 1.304, 
    1.294, 1.281, 1.266, 1.251, 1.235, 1.219, 1.203, 1.186, 1.169, 1.151, 
    1.133, 1.115, 1.097, 1.079, 1.062, 1.046, 1.031, 1.019, 1.009, 1.003, 
    0.999, 0.999, 1.001, 1.004, 1.007, 1.009, 1.008, 1.004, 0.999, 0.993, 
    0.992, 0.998, 1.018, 1.055, 1.109, 1.175, 1.247, 1.314, 1.383, 1.486, 
    1.674, 1.942, 2.143, 2.168, 2.08, 1.954, 1.817, 1.678, 1.538, 1.407, 
    1.315, 1.314, 1.451, 1.721, 2.019, 2.328, 2.744, 3.046, 3.073, 2.968, 
    2.843, 2.73, 2.634, 2.554, 2.486, 2.428, 2.379, 2.335, 2.297, 2.263, 
    2.233, 2.206, 2.181, 2.158 ;

 idx_rfr_montmorillonite_img = 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.005, 0.005, 0.005, 0.006, 
    0.007, 0.008, 0.01, 0.013, 0.019, 0.028, 0.033, 0.025, 0.017, 0.012, 
    0.009, 0.008, 0.007, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 
    0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 
    0.006, 0.006, 0.006, 0.006, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 
    0.007, 0.007, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.01, 0.01, 0.01, 0.01, 0.01, 0.011, 0.011, 
    0.011, 0.011, 0.012, 0.012, 0.012, 0.013, 0.013, 0.013, 0.014, 0.014, 
    0.014, 0.015, 0.015, 0.015, 0.016, 0.016, 0.017, 0.017, 0.018, 0.018, 
    0.019, 0.02, 0.02, 0.021, 0.022, 0.023, 0.023, 0.024, 0.025, 0.026, 
    0.027, 0.028, 0.029, 0.031, 0.032, 0.034, 0.035, 0.037, 0.039, 0.041, 
    0.043, 0.045, 0.048, 0.05, 0.053, 0.057, 0.061, 0.065, 0.07, 0.075, 
    0.081, 0.088, 0.096, 0.105, 0.116, 0.129, 0.144, 0.163, 0.185, 0.212, 
    0.244, 0.282, 0.326, 0.375, 0.426, 0.478, 0.53, 0.582, 0.636, 0.691, 
    0.742, 0.78, 0.793, 0.774, 0.737, 0.706, 0.697, 0.718, 0.768, 0.841, 
    0.931, 1.03, 1.14, 1.25, 1.37, 1.49, 1.62, 1.74, 1.84, 1.9, 1.89, 1.82, 
    1.68, 1.54, 1.43, 1.37, 1.31, 1.22, 1.08, 0.919, 0.759, 0.623, 0.514, 
    0.43, 0.364, 0.313, 0.272, 0.24, 0.214, 0.193, 0.176, 0.162, 0.151, 
    0.142, 0.136, 0.132, 0.13, 0.133, 0.139, 0.152, 0.174, 0.204, 0.234, 
    0.242, 0.218, 0.183, 0.155, 0.136, 0.128, 0.128, 0.135, 0.145, 0.15, 
    0.141, 0.123, 0.106, 0.093, 0.086, 0.086, 0.093, 0.099, 0.086, 0.07, 
    0.06, 0.054, 0.051, 0.05, 0.049, 0.05, 0.051, 0.054, 0.059, 0.067, 0.078, 
    0.092, 0.097, 0.089, 0.075, 0.064, 0.057, 0.052, 0.05, 0.048, 0.047, 
    0.047, 0.047, 0.048, 0.049, 0.05, 0.051, 0.053, 0.055, 0.057, 0.06, 
    0.064, 0.068, 0.075, 0.083, 0.092, 0.093, 0.091, 0.092, 0.095, 0.1, 
    0.106, 0.113, 0.122, 0.131, 0.142, 0.155, 0.169, 0.186, 0.204, 0.225, 
    0.248, 0.274, 0.303, 0.334, 0.367, 0.401, 0.436, 0.47, 0.503, 0.535, 
    0.564, 0.594, 0.624, 0.657, 0.696, 0.743, 0.8, 0.866, 0.94, 1.02, 1.09, 
    1.15, 1.2, 1.24, 1.3, 1.38, 1.45, 1.4, 1.18, 0.921, 0.731, 0.621, 0.572, 
    0.572, 0.624, 0.739, 0.932, 1.19, 1.47, 1.66, 1.72, 1.75, 1.64, 1.27, 
    0.864, 0.592, 0.425, 0.321, 0.253, 0.206, 0.172, 0.147, 0.127, 0.112, 
    0.099, 0.089, 0.081, 0.073, 0.067, 0.062 ;
}

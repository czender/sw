// ncgen -b -o ~ammann/DATA/AERO/idx_rfr/idx_rfr_PaW75.nc ~ammann/DATA/AERO/idx_rfr/idx_rfr_PaW75.cdl
// ncks -C -H -s %9.5f -v bnd,idx_rfr_H2SO4_300K_PaW75_img,idx_rfr_H2SO4_300K_PaW75_rl /ammann/DATA/AERO/idx_rfr/idx_rfr_PaW75.nc

netcdf idx_rfr_PaW75 {
dimensions:
        bnd=236;
        bnd_HSL88=62;
variables:
        :history = "";
        :source="Thu Jun 20 MDT 1999
PaW75 : from palmer_w.dat in $HOME/idx_rfr/hitran
PaW75 : Kent F. Palmer and Dudley Williams, 1975: Optical constants of sulfuric acid; application to the clouds of Venus? Applied Optics 14, 1, p. 208-219.
PaW75 : Range 0.36--25.0 microns; extended 0.33-0.2 and 27-50 micron with HSL88. These indices are also shown graphically in PaW75.
PaW75 : File in HITRAN provides values at 25%, 38%, 50%, 75%, 84.5%, 95.6% H2SO4 solutions (by weight)
PaW75 : Values below are for 75% H2SO4 (and 25% H2O) by weight
HSL88 : from /home/zender/idx_rfr/hitran/shettle.dat
HSL88 : Hummel, J. R., Shettle, E. P. and Longtin, D. R. (1988) A New Background Stratospheric Aerosol Model for Use in Atmospheric Radiation Models, AFGL-TR-88-0166, Air Force Geophysics Laboratory, Hanscom AFB, MA, August 1988.
HSL88 : Range used : 0.2 - 0.337 micron, optical constants for H2SO4 75% for 300 (here only 300K).";

        float bnd(bnd);
        bnd:long_name = "Band center wavelength";
        bnd:units = "micron";
        bnd:C_format = "%.3g";

        float bnd_HSL88(bnd_HSL88);
        bnd_HSL88:long_name = "Band center wavelength";
        bnd_HSL88:units = "micron";
        bnd_HSL88:C_format = "%.5g";

        float idx_rfr_H2SO4_300K_PaW75_rl(bnd);
        idx_rfr_H2SO4_300K_PaW75_rl:long_name = "Sulfate 75% real index of refraction";
        idx_rfr_H2SO4_300K_PaW75_rl:units = "";
        idx_rfr_H2SO4_300K_PaW75_rl:C_format = "%.3g";

        float idx_rfr_H2SO4_300K_PaW75_img(bnd);
        idx_rfr_H2SO4_300K_PaW75_img:long_name = "Sulfate 75% imaginary index of refraction";
        idx_rfr_H2SO4_300K_PaW75_img:units = "";
        idx_rfr_H2SO4_300K_PaW75_img:C_format = "%.5g";

        float idx_rfr_H2SO4_300K_75_HSL88_rl(bnd_HSL88);
        idx_rfr_H2SO4_300K_75_HSL88_rl:long_name = "Sulfate 75% real index of refraction";
        idx_rfr_H2SO4_300K_75_HSL88_rl:units = "";
        idx_rfr_H2SO4_300K_75_HSL88_rl:C_format = "%.3g";

        float idx_rfr_H2SO4_300K_75_HSL88_img(bnd_HSL88);
        idx_rfr_H2SO4_300K_75_HSL88_img:long_name = "Sulfate 75% imaginary index of refraction";
        idx_rfr_H2SO4_300K_75_HSL88_img:units = "";
        idx_rfr_H2SO4_300K_75_HSL88_img:C_format = "%.5g";


data:


bnd =
 50.000, 40.000, 35.000, 30.000, 27.900, 
 25.000, 24.390, 23.256, 22.727, 22.222, 21.277, 20.833, 20.408, 20.000, 19.608, 18.868, 18.519, 18.182, 17.857, 17.544, 17.241, 16.949, 16.667, 16.129, 15.873, 15.385, 14.925, 14.706, 14.286, 13.889, 13.514, 13.158, 12.821, 12.658, 12.500, 12.195, 11.905, 11.765, 11.494, 11.442, 11.364, 11.236, 11.111, 10.989, 10.870, 10.753, 10.638, 10.526, 10.417, 10.384, 10.309, 10.204, 10.101,  9.901,  9.804,  9.709,  9.615,  9.524,  9.434,  9.346,  9.259,  9.174,  9.091,  9.009,  8.929,  8.850,  8.696,  8.621,  8.547,  8.403,  8.264,  8.130,  8.065,  8.000,  7.874,  7.752,  7.634,  7.576,  7.463,  7.353,  7.299,  7.194,  7.092,  6.993,  6.897,  6.803,  6.711,  6.667,  6.623,  6.579,  6.536,  6.494,  6.410,  6.329,  6.250,  6.211,  6.173,  6.135,  6.098,  6.061,  6.024,  5.952,  5.882,  5.814,  5.747,  5.682,  5.650,  5.618,  5.556,  5.495,  5.435,  5.376,  5.319,  5.263,  5.181,  5.102,  4.950,  4.808,  4.717,  4.587,  4.464,  4.367,  4.292,  4.274,  4.219,  4.149,  4.082,  4.000,  3.953,  3.906,  3.861,  3.846,  3.817,  3.759,  3.690,  3.623,  3.559,  3.472,  3.413,  3.344,  3.279,  3.175,  3.077,  3.021,  2.985,  2.941,  2.915,  2.882,  2.841,  2.833,  2.770,  2.762,  2.725,  2.688,  2.632,  2.564,  2.500,  2.439,  2.381,  2.326,  2.273,  2.222,  2.174,  2.128,  2.083,  2.041,  2.000,  1.961,  1.923,  1.887,  1.852,  1.818,  1.786,  1.754,  1.724,  1.695,  1.667,  1.639,  1.613,  1.587,  1.562,  1.538,  1.515,  1.493,  1.471,  1.449,  1.429,  1.408,  1.389,  1.370,  1.351,  1.333,  1.316,  1.299,  1.282,  1.266,  1.250,  1.220,  1.190,  1.163,  1.136,  1.111,  1.087,  1.064,  1.042,  1.020,  1.000,   .980,   .962,   .943,   .926,   .909,   .893,   .877,   .862,   .847,   .833,   .820,   .806,   .794,   .781,   .769,   .758,   .746,   .735,   .725,   .714,   .702,   .556,   .449,   .445,   .360,
 .337,   .300,   .250,   .200  ;


 idx_rfr_H2SO4_300K_PaW75_rl =
 2.010, 1.940, 1.720, 1.730, 1.780,
 1.930, 1.939, 1.918, 1.881, 1.848, 1.781, 1.782, 1.804, 1.823, 1.842, 1.892, 1.926, 1.946, 1.939, 1.869, 1.741, 1.621, 1.542, 1.512, 1.512, 1.551, 1.596, 1.613, 1.643, 1.663, 1.681, 1.701, 1.726, 1.741, 1.757, 1.796, 1.844, 1.869, 1.916, 1.911, 1.904, 1.842, 1.739, 1.676, 1.663, 1.678, 1.717, 1.756, 1.788, 1.807, 1.822, 1.849, 1.882, 1.947, 1.944, 1.907, 1.807, 1.702, 1.624, 1.589, 1.590, 1.626, 1.655, 1.669, 1.666, 1.643, 1.545, 1.479, 1.421, 1.320, 1.241, 1.179, 1.161, 1.151, 1.145, 1.144, 1.136, 1.133, 1.142, 1.173, 1.192, 1.222, 1.249, 1.272, 1.297, 1.308, 1.323, 1.331, 1.340, 1.351, 1.361, 1.368, 1.384, 1.399, 1.413, 1.422, 1.428, 1.434, 1.433, 1.430, 1.427, 1.420, 1.410, 1.392, 1.371, 1.361, 1.356, 1.350, 1.341, 1.337, 1.336, 1.336, 1.339, 1.342, 1.347, 1.353, 1.366, 1.379, 1.384, 1.386, 1.384, 1.386, 1.395, 1.397, 1.405, 1.399, 1.400, 1.398, 1.396, 1.395, 1.395, 1.395, 1.396, 1.396, 1.397, 1.394, 1.388, 1.370, 1.357, 1.341, 1.325, 1.306, 1.296, 1.294, 1.292, 1.288, 1.284, 1.277, 1.273, 1.272, 1.277, 1.279, 1.293, 1.308, 1.320, 1.332, 1.344, 1.352, 1.358, 1.362, 1.367, 1.370, 1.374, 1.377, 1.380, 1.382, 1.384, 1.386, 1.388, 1.389, 1.391, 1.392, 1.393, 1.394, 1.396, 1.397, 1.398, 1.398, 1.399, 1.400, 1.402, 1.403, 1.403, 1.404, 1.405, 1.406, 1.406, 1.407, 1.408, 1.409, 1.410, 1.410, 1.411, 1.411, 1.412, 1.413, 1.413, 1.415, 1.416, 1.416, 1.417, 1.418, 1.419, 1.420, 1.421, 1.421, 1.422, 1.422, 1.423, 1.423, 1.424, 1.424, 1.425, 1.425, 1.425, 1.426, 1.426, 1.427, 1.427, 1.427, 1.427, 1.427, 1.427, 1.427, 1.427, 1.427, 1.427, 1.428, 1.431, 1.432, 1.438, 1.452,
1.459, 1.469, 1.484, 1.498  ;


 idx_rfr_H2SO4_300K_PaW75_img =
 0.650, 0.630, 0.520, 0.290, 0.250,
 2.00E-01, 2.26E-01, 3.00E-01, 3.20E-01, 3.29E-01, 2.90E-01, 2.57E-01, 2.40E-01, 2.35E-01, 2.38E-01, 2.61E-01, 2.99E-01, 3.62E-01, 4.57E-01, 5.54E-01, 5.94E-01, 5.64E-01, 4.79E-01, 3.52E-01, 2.99E-01, 2.21E-01, 1.91E-01, 1.83E-01, 1.73E-01, 1.71E-01, 1.65E-01, 1.60E-01, 1.57E-01, 1.57E-01, 1.58E-01, 1.68E-01, 1.94E-01, 2.16E-01, 3.13E-01, 3.41E-01, 3.86E-01, 4.64E-01, 4.63E-01, 4.10E-01, 3.51E-01, 3.01E-01, 2.75E-01, 2.71E-01, 2.77E-01, 2.82E-01, 2.92E-01, 3.11E-01, 3.38E-01, 4.53E-01, 5.38E-01, 6.37E-01, 7.08E-01, 7.11E-01, 6.68E-01, 6.12E-01, 5.60E-01, 5.40E-01, 5.56E-01, 5.90E-01, 6.34E-01, 6.81E-01, 7.55E-01, 7.61E-01, 7.58E-01, 7.19E-01, 6.63E-01, 5.93E-01, 5.47E-01, 5.13E-01, 4.45E-01, 3.97E-01, 3.51E-01, 3.23E-01, 2.62E-01, 2.11E-01, 1.95E-01, 1.73E-01, 1.58E-01, 1.43E-01, 1.43E-01, 1.37E-01, 1.30E-01, 1.26E-01, 1.22E-01, 1.21E-01, 1.22E-01, 1.23E-01, 1.25E-01, 1.30E-01, 1.38E-01, 1.44E-01, 1.52E-01, 1.64E-01, 1.75E-01, 1.84E-01, 1.91E-01, 2.03E-01, 2.15E-01, 2.25E-01, 2.20E-01, 2.12E-01, 2.09E-01, 2.06E-01, 1.94E-01, 1.82E-01, 1.71E-01, 1.60E-01, 1.51E-01, 1.44E-01, 1.35E-01, 1.28E-01, 1.18E-01, 1.16E-01, 1.17E-01, 1.21E-01, 1.19E-01, 1.13E-01, 1.09E-01, 1.10E-01, 1.17E-01, 1.21E-01, 1.24E-01, 1.26E-01, 1.27E-01, 1.27E-01, 1.27E-01, 1.27E-01, 1.28E-01, 1.30E-01, 1.36E-01, 1.43E-01, 1.53E-01, 1.61E-01, 1.59E-01, 1.59E-01, 1.50E-01, 1.31E-01, 1.09E-01, 9.90E-02, 9.30E-02, 8.60E-02, 8.20E-02, 7.30E-02, 5.60E-02, 5.20E-02, 2.30E-02, 1.90E-02, 6.00E-03, 0.00E+00, 0.00E+00, 0.00E+00, 3.76E-03, 2.97E-03, 2.41E-03, 2.09E-03, 1.86E-03, 1.67E-03, 1.54E-03, 1.43E-03, 1.35E-03, 1.30E-03, 1.26E-03, 1.24E-03, 1.11E-03, 7.96E-04, 5.95E-04, 5.37E-04, 4.86E-04, 4.24E-04, 3.61E-04, 3.14E-04, 2.72E-04, 2.34E-04, 2.02E-04, 1.76E-04, 1.55E-04, 1.38E-04, 1.25E-04, 1.17E-04, 1.10E-04, 1.02E-04, 8.78E-05, 6.16E-05, 3.89E-05, 2.59E-05, 1.98E-05, 1.59E-05, 1.27E-05, 1.05E-05, 8.93E-06, 7.75E-06, 6.94E-06, 5.63E-06, 4.95E-06, 4.05E-06, 2.46E-06, 1.84E-06, 1.60E-06, 1.50E-06, 1.48E-06, 1.52E-06, 1.53E-06, 1.41E-06, 1.03E-06, 6.05E-07, 3.62E-07, 2.84E-07, 2.33E-07, 2.02E-07, 1.83E-07, 1.58E-07, 1.24E-07, 9.98E-08, 8.79E-08, 8.46E-08, 8.39E-08, 8.20E-08, 7.84E-08, 6.83E-08, 4.80E-08, 3.58E-08, 2.79E-08, 2.07E-08, 0.00E+00, 0.00E+00, 0.00E+00, 0.00E+00,  
 1.00E-8, 1.00E-8, 1.00E-8, 1.00E-8  ;

 bnd_HSL88 =
 0.200, 0.250, 0.300, 0.337, 0.400, 0.488, 0.515, 0.550, 0.633, 0.694, 0.860, 1.060, 1.300, 1.536, 1.800, 2.000, 2.250, 2.500, 2.700, 3.000, 3.200, 3.392, 3.500, 3.750, 4.000, 4.500, 5.000, 5.500, 6.000, 6.200, 6.500, 7.200, 7.900, 8.200, 8.500, 8.700, 9.000, 9.200, 9.500, 9.800,  10.000,  10.591,  11.000,  11.500,  12.500,  13.000,  14.000,  14.800,  15.000,  16.400,  17.200,  18.000,  18.500,  20.000,  21.300,  22.500,  25.000,  27.900,  30.000,  35.000,  40.000,  50.000  ;

 idx_rfr_H2SO4_300K_75_HSL88_rl =
 1.498, 1.484, 1.469, 1.459, 1.440, 1.432, 1.431, 1.430, 1.429, 1.428, 1.425, 1.420, 1.410, 1.403, 1.390, 1.384, 1.370, 1.344, 1.303, 1.293, 1.311, 1.352, 1.376, 1.396, 1.398, 1.385, 1.360, 1.337, 1.425, 1.424, 1.370, 1.210, 1.140, 1.200, 1.370, 1.530, 1.650, 1.600, 1.670, 1.910, 1.890, 1.720, 1.670, 1.890, 1.740, 1.690, 1.640, 1.610, 1.590, 1.520, 1.724, 1.950, 1.927, 1.810, 1.790, 1.820, 1.840, 1.780, 1.730, 1.720, 1.940, 2.010  ;

 idx_rfr_H2SO4_300K_75_HSL88_img =
 1.00E-8, 1.00E-8, 1.00E-8, 1.00E-8, 1.00E-8, 1.00E-8, 1.00E-8, 1.00E-8, 1.47E-8, 1.99E-8, 1.79E-7, 1.50E-6, 1.00E-5, 1.37E-4, 5.50E-4, 0.00126, 0.00180, 0.00376, 0.00570, 0.0955, 0.135, 0.159, 0.158, 0.131, 0.126, 0.120, 0.121, 0.183, 0.195, 0.165, 0.128, 0.176, 0.488, 0.645, 0.755, 0.772, 0.633, 0.586, 0.750, 0.680, 0.455, 0.340, 0.485, 0.374, 0.198, 0.195, 0.195, 0.205, 0.211, 0.414, 0.590, 0.410, 0.302, 0.230, 0.250, 0.290, 0.240, 0.250, 0.290, 0.520, 0.630, 0.650  ;


}

























// $Id$
// ncgen -b -o ${DATA}/aca/idx_rfr_shettle.nc ${HOME}/idx_rfr/idx_rfr_shettle.cdl

netcdf idx_rfr_shettle {
dimensions:
	bnd=62;
variables:

	:RCS_Header = "$Id$";
	:history = "";
	:source="HITRAN96 CDROM file /cdrom/aerosols/shettle.dat,
Table A4";

	float bnd(bnd);
	bnd:long_name = "Band center wavelength";
	bnd:units = "micron";
	bnd:C_format = "%.5g";

	float idx_rfr_h2so4_215K_rl(bnd);
	idx_rfr_h2so4_215K_rl:long_name = "75% H2SO4 25% H2O (by weight) at 215K real index of refraction";
	idx_rfr_h2so4_215K_rl:units = "";
	idx_rfr_h2so4_215K_rl:composition = "75% H2SO4 25% H2O (by weight)";
	idx_rfr_h2so4_215K_rl:C_format = "%.4g";

	float idx_rfr_h2so4_215K_img(bnd);
	idx_rfr_h2so4_215K_img:long_name = "75% H2SO4 25% H2O (by weight) at 215K imaginary index of refraction";
	idx_rfr_h2so4_215K_img:units = "";
	idx_rfr_h2so4_215K_img:composition = "75% H2SO4 25% H2O (by weight)";
	idx_rfr_h2so4_215K_img:C_format = "%.3g";

	float idx_rfr_h2so4_300K_rl(bnd);
	idx_rfr_h2so4_300K_rl:long_name = "75% H2SO4 25% H2O (by weight) at 300K real index of refraction";
	idx_rfr_h2so4_300K_rl:units = "";
	idx_rfr_h2so4_300K_rl:composition = "75% H2SO4 25% H2O (by weight)";
	idx_rfr_h2so4_300K_rl:C_format = "%.4g";

	float idx_rfr_h2so4_300K_img(bnd);
	idx_rfr_h2so4_300K_img:long_name = "75% H2SO4 25% H2O (by weight) at 300K imaginary index of refraction";
	idx_rfr_h2so4_300K_img:units = "";
	idx_rfr_h2so4_300K_img:composition = "75% H2SO4 25% H2O (by weight)";
	idx_rfr_h2so4_300K_img:C_format = "%.3g";

	float idx_rfr_volcanic_dust_rl(bnd);
	idx_rfr_volcanic_dust_rl:long_name = "Volcanic dust real index of refraction";
	idx_rfr_volcanic_dust_rl:units = "";
	idx_rfr_volcanic_dust_rl:C_format = "%.4g";

	float idx_rfr_volcanic_dust_img(bnd);
	idx_rfr_volcanic_dust_img:long_name = "Volcanic dust imaginary index of refraction";
	idx_rfr_volcanic_dust_img:units = "";
	idx_rfr_volcanic_dust_img:C_format = "%.3g";

	float idx_rfr_meteoric_dust_rl(bnd);
	idx_rfr_meteoric_dust_rl:long_name = "Meteoric dust real index of refraction";
	idx_rfr_meteoric_dust_rl:units = "";
	idx_rfr_meteoric_dust_rl:C_format = "%.4g";

	float idx_rfr_meteoric_dust_img(bnd);
	idx_rfr_meteoric_dust_img:long_name = "Meteoric dust imaginary index of refraction";
	idx_rfr_meteoric_dust_img:units = "";
	idx_rfr_meteoric_dust_img:C_format = "%.3g";

data:	
 bnd = 0.200,  0.250,  0.300,  0.337,  0.400,  0.488,  0.515,  0.550,
	0.633, 	0.694,  0.860,  1.060,  1.300,  1.536,  1.800,  2.000,
	2.250, 	2.500,  2.700, 	3.000,  3.200,  3.392,  3.500,  3.750,
	4.000, 	4.500,  5.000,  5.500,  6.000, 	6.200,  6.500,  7.200,
	7.900,  8.200,  8.500,  8.700,  9.000,  9.200,  9.500,  9.800,
	10.000, 10.591, 11.000, 11.500, 12.500, 13.000, 14.000, 14.800,  
	15.000, 16.400, 17.200, 18.000, 18.500, 20.000, 21.300, 22.500,
	25.000, 27.900, 30.000, 35.000, 40.000, 50.000;  
 
 idx_rfr_volcanic_dust_rl = 
	1.500, 1.500, 1.500, 1.500, 1.500, 1.500, 1.500, 1.500, 1.500, 1.500,
	1.500, 1.500, 1.500, 1.490, 1.480, 1.460, 1.460, 1.460, 1.460, 1.480,
	1.480, 1.490, 1.490, 1.500, 1.500, 1.520, 1.510, 1.510, 1.480, 1.460,
	1.450, 1.440, 1.380, 1.340, 1.620, 1.950, 2.200, 2.230, 2.250, 2.280,
	2.300, 2.200, 2.150, 2.050, 1.800, 1.760, 1.700, 1.650, 1.650, 1.750,
	1.850, 2.000, 2.100, 2.250, 2.400, 2.500, 2.600, 2.500, 2.400, 2.300,
	2.250, 0.000; 
 idx_rfr_volcanic_dust_img = 
	0.070, 0.030, 0.010, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008,
	0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.009, 0.010, 0.013,
	0.014, 0.012, 0.011, 0.009, 0.007, 0.0075, 0.0090, 0.012, 0.015,
	0.018, 0.024, 0.045, 0.072, 0.097, 0.121, 0.170, 0.215, 0.240, 0.275,
	0.304, 0.320, 0.305, 0.270, 0.240, 0.155, 0.148, 0.145, 0.157, 0.170,
	0.200, 0.240, 0.305, 0.325, 0.318, 0.290, 0.350, 0.400, 0.430, 0.450,
	0.520, 0.650, 0.000;

 idx_rfr_h2so4_215K_rl = 
	1.526, 1.512, 1.496, 1.484, 1.464, 1.456, 1.454, 1.454, 1.452, 1.452,
	1.448, 1.443, 1.432, 1.425, 1.411, 1.405, 1.390, 1.362, 1.319, 1.288,
	1.292, 1.366, 1.383, 1.420, 1.435, 1.427, 1.411, 1.376, 1.485, 1.485,
	1.421, 1.235, 1.148, 1.220, 1.457, 1.753, 1.767, 1.704, 1.791, 2.128,
	2.094, 1.805, 1.823, 2.024, 1.808, 1.790, 1.739, 1.663, 1.656, 1.692,
	2.003, 2.207, 2.041, 1.895, 1.809, 1.942, 1.993, 0.000, 0.000, 0.000,
	0.000, 0.000;
 idx_rfr_h2so4_215K_img = 
	1.07e-8, 1.07e-8, 1.07e-8, 1.07e-8, 1.07e-8, 1.07e-8, 1.07e-8,
	1.07e-8, 1.56e-8, 2.12e-8, 1.90e-7, 1.60e-6, 1.06e-5, 1.46e-4,
	5.85e-4, 0.00134, 0.00192, 0.00399, 0.00604, 0.0875, 0.144, 0.178,
	0.179, 0.165, 0.151, 0.156, 0.137, 0.195, 0.195, 0.147,
	0.0841, 0.166, 0.461, 0.709, 0.840, 0.817, 0.604, 0.557,
	0.736, 0.465, 0.306, 0.210, 0.433, 0.199, 0.110, 0.112,
	0.134, 0.163, 0.181, 0.463, 0.616, 0.166, 0.0940,
	0.0558, 0.146, 0.187, 0.0274, 0.000, 0.000, 0.000, 0.000,
	0.000;  

 idx_rfr_h2so4_300K_rl = 
	1.498, 1.484, 1.469, 1.459, 1.440, 1.432, 1.431, 1.430, 1.429, 1.428,
	1.425, 1.420, 1.410, 1.403, 1.390, 1.384, 1.370, 1.344, 1.303, 1.293,
	1.311, 1.352, 1.376, 1.396, 1.398, 1.385, 1.360, 1.337, 1.425, 1.424,
	1.370, 1.210, 1.140, 1.200, 1.370, 1.530, 1.650, 1.600, 1.670, 1.910,
	1.890, 1.720, 1.670, 1.890, 1.740, 1.690, 1.640, 1.610, 1.590, 1.520,
	1.724, 1.950, 1.927, 1.810, 1.790, 1.820, 1.840, 1.780, 1.730, 1.720,
	1.940, 2.010; 
 idx_rfr_h2so4_300K_img = 
	1.00e-8, 1.00e-8, 1.00e-8, 1.00e-8, 1.00e-8, 1.00e-8, 1.00e-8,
	1.00e-8, 1.47e-8, 1.99e-8, 1.79e-7, 1.50e-6, 1.00e-5, 1.37e-4,
	5.50e-4, 0.00126, 0.00180, 0.00376, 0.00570, 0.0955, 0.135, 0.159,
	0.158, 0.131, 0.126, 0.120, 0.121, 0.183, 0.195, 0.165,
	0.128, 0.176, 0.488, 0.645, 0.755, 0.772, 0.633, 0.586,
	0.750, 0.680, 0.455, 0.340, 0.485, 0.374, 0.198, 0.195,
	0.195, 0.205, 0.211, 0.414, 0.590, 0.410, 0.302, 0.230,
	0.250, 0.290, 0.240, 0.250, 0.290, 0.520, 0.630, 0.650;  

 idx_rfr_meteoric_dust_rl = 
	1.515, 1.515, 1.515, 1.514, 1.514, 1.513, 1.513, 1.513, 1.512, 1.511,
	1.509, 1.506, 1.501, 1.495, 1.488, 1.482, 1.474, 1.467, 1.462, 1.456,
	1.454, 1.454, 1.455, 1.459, 1.466, 1.485, 1.500, 1.508, 1.507, 1.504,
	1.497, 1.469, 1.422, 1.395, 1.363, 1.339, 1.302, 1.281, 1.272, 1.310,
	1.355, 1.419, 1.509, 1.847, 1.796, 1.711, 1.641, 1.541, 1.510, 1.478,
	1.441, 1.354, 1.389, 1.803, 1.797, 1.661, 1.983, 2.023, 2.149, 2.146,
	1.979, 0.000; 
 idx_rfr_meteoric_dust_img = 
	1.23e-5, 2.41e-5, 4.18e-5, 5.94e-5, 9.95e-5, 1.81e-4, 2.13e-4,
	2.61e-4, 3.99e-4, 5.30e-4, 0.00102, 0.00195, 0.00372, 0.00634, 0.0106,
	0.0151, 0.0224, 0.0318, 0.0410, 0.0573, 0.0694, 0.0815,
	0.0882, 0.103, 0.116, 0.131, 0.135, 0.132, 0.126, 0.124,
	0.121, 0.119, 0.130, 0.142, 0.162, 0.182, 0.228, 0.273,
	0.360, 0.450, 0.488, 0.547, 0.691, 0.634, 0.252, 0.219,
	0.217, 0.198, 0.206, 0.467, 0.400, 0.557, 0.705, 0.765,
	0.556, 0.592, 0.861, 0.666, 0.665, 0.380, 0.359, 0.000;  
}

// ncgen -b -o ${DATA}/aca/idx_rfr_Vol73.nc ${HOME}/idx_rfr/idx_rfr_Vol73.cdl
// ncks -C -H -d bnd,0.5e-6 -v idx_rfr_saharan_dust_img,idx_rfr_saharan_dust_rl ${DATA}/aca/idx_rfr_Vol73.nc

netcdf idx_rfr_Vol73 {

dimensions:
	bnd_Pat81=23;
	bnd_Vol73=1993;
	bnd=2023;
variables:

	:RCS_Header = "$Id$";
	:history = "";
	:source="
Tue Jun  9 15:08:40 MDT 1998:
Added saharan_dust, which is a combination of Pat81, DKS91, and Vol73. 
Pat81 and Vol73 optical properties were supplied by Irina Sokolik.
Pat81 data are 23 measurements of n+ik between 0.25005 and 0.69005 microns.
Vol73 data are 1993 measurements of n+ik between 2.5813 and 39.084 microns.
saharan_dust uses afghan_dust to fill in the gaps in the SW.
afghan dust data are used for 6 bands from 0.71429--2.564 microns.
The afghan_dust data come from SAJ93, as stored in ${HOME}/dst/idx_rfr_SAJ93.nc.
mineral_dust data are used for the band at 0.2 microns.
The mineral_dust data come from DKS91, as stored in ${HOME}/dst/idx_rfr_dks91.nc.
Saharan dust is much more optically active than dust_like or mineral_dust aerosols of DKS91.";

	float bnd(bnd);
	bnd:long_name = "Band center wavelength";
	bnd:units = "micron";
	bnd:C_format = "%.5g";

	float bnd_Pat81(bnd_Pat81);
	bnd_Pat81:long_name = "Band center wavelength";
	bnd_Pat81:units = "micron";
	bnd_Pat81:C_format = "%.5g";

	float bnd_Vol73(bnd_Vol73);
	bnd_Vol73:long_name = "Band center wavelength";
	bnd_Vol73:units = "micron";
	bnd_Vol73:C_format = "%.5g";

	float idx_rfr_saharan_dust_rl(bnd);
	idx_rfr_saharan_dust_rl:long_name = "Saharan dust real index of refraction";
	idx_rfr_saharan_dust_rl:units = "";
	idx_rfr_saharan_dust_rl:C_format = "%.4g";

	float idx_rfr_saharan_dust_img(bnd);
	idx_rfr_saharan_dust_img:long_name = "Saharan dust imaginary index of refraction";
	idx_rfr_saharan_dust_img:units = "";
	idx_rfr_saharan_dust_img:C_format = "%.3g";

	float idx_rfr_Pat81_rl(bnd_Pat81);
	idx_rfr_Pat81_rl:long_name = "Saharan dust real index of refraction";
	idx_rfr_Pat81_rl:units = "";
	idx_rfr_Pat81_rl:C_format = "%.4g";

	float idx_rfr_Pat81_img(bnd_Pat81);
	idx_rfr_Pat81_img:long_name = "Saharan dust imaginary index of refraction";
	idx_rfr_Pat81_img:units = "";
	idx_rfr_Pat81_img:C_format = "%.3g";

	float idx_rfr_Vol73_rl(bnd_Vol73);
	idx_rfr_Vol73_rl:long_name = "Saharan dust real index of refraction";
	idx_rfr_Vol73_rl:units = "";
	idx_rfr_Vol73_rl:C_format = "%.4g";

	float idx_rfr_Vol73_img(bnd_Vol73);
	idx_rfr_Vol73_img:long_name = "Saharan dust imaginary index of refraction";
	idx_rfr_Vol73_img:units = "";
	idx_rfr_Vol73_img:C_format = "%.3g";

data:	

bnd_Pat81 = 0.2500,0.2700,0.2900,0.3100,0.3300,0.3500,0.3700,0.3900,0.4100,0.4300,0.4500,0.4700,0.4900,0.5100,0.5300,0.5500,0.5700,0.5900,0.6100,0.6300,0.6500,0.6700,0.6900;
idx_rfr_Pat81_rl = 1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56;
idx_rfr_Pat81_img = 0.050561,0.045743,0.038785,0.031728,0.027208,0.023094,0.019765,0.016975,0.014397,0.012447,0.010859,0.009481,0.008340,0.007342,0.006425,0.005638,0.004929,0.004435,0.003992,0.003811,0.003810,0.003774,0.003773;

bnd = 0.2, 
0.2500,0.2700,0.2900,0.3100,0.3300,0.3500,0.3700,0.3900,0.4100,0.4300,0.4500,0.4700,0.4900,0.5100,0.5300,0.5500,0.5700,0.5900,0.6100,0.6300,0.6500,0.6700,0.6900,
0.714290,0.769230,0.833330,0.909090,2.500000,2.564100,
2.5813,2.5995,2.6178,2.63605,2.65431,2.67256,2.69081,2.70906,2.72731,2.74556,2.76381,2.78206,2.80032,2.8185,2.83682,2.85507,2.87332,2.89157,2.90982,2.92808,2.94633,2.96458,2.98283,3.00108,3.01933,3.03758,3.05584,3.07409,3.09234,3.11059,3.12884,3.14709,3.16534,3.18359,3.20185,3.2201,3.23835,3.2566,3.27485,3.2931,3.31135,3.32961,3.34786,3.36611,3.38436,3.40261,3.42086,3.43911,3.45736,3.47562,3.49387,3.51212,3.53037,3.54862,3.56687,3.58512,3.60338,3.62163,3.63988,3.65813,3.67638,3.69463,3.71288,3.73114,3.74939,3.76764,3.78589,3.80414,3.82239,3.84064,3.85889,3.87715,3.8954,3.91365,3.9319,3.95015,3.9684,3.98665,4.00491,4.02316,4.04141,4.05966,4.07791,4.09616,4.11441,4.13266,4.15092,4.16917,4.18742,4.20567,4.22392,4.24217,4.26042,4.27868,4.29693,4.31518,4.33343,4.35168,4.36993,4.38818,4.40643,4.42469,4.44294,4.46119,4.47944,4.49769,4.51594,4.53419,4.55245,4.5707,4.58895,4.6072,4.62545,4.6437,4.66195,4.68021,4.69846,4.71671,4.73496,4.75321,4.77146,4.78971,4.80796,4.82622,4.84447,4.86272,4.88097,4.89922,4.91747,4.93572,4.95398,4.97223,4.99048,5.00873,5.02698,5.04523,5.06348,5.08173,5.09999,5.11824,5.13649,5.15474,5.17299,5.19124,5.20949,5.22775,5.246,5.26425,5.2825,5.30075,5.319,5.33725,5.35551,5.37376,5.39201,5.41026,5.42851,5.44676,5.46501,5.48326,5.50152,5.51977,5.53802,5.55627,5.57452,5.59277,5.61102,5.62928,5.64753,5.66578,5.68403,5.70228,5.72053,5.73878,5.75703,5.77529,5.79354,5.81179,5.83004,5.84829,5.86654,5.88479,5.90305,5.9213,5.93955,5.9578,5.97605,5.9943,6.01255,6.03081,6.04906,6.06731,6.08556,6.10381,6.12206,6.14031,6.15856,6.17682,6.19507,6.21332,6.23157,6.24982,6.26807,6.28632,6.30458,6.32283,6.34108,6.35933,6.37758,6.39583,6.41408,6.43233,6.45059,6.46884,6.48709,6.50534,6.52359,6.54184,6.56009,6.57835,6.5966,6.61485,6.6331,6.65135,6.6696,6.68785,6.70611,6.72436,6.74261,6.76086,6.77911,6.79736,6.81561,6.83386,6.85212,6.87037,6.88862,6.90687,6.92512,6.94337,6.96162,6.97988,6.99813,7.01638,7.03463,7.05288,7.07113,7.08938,7.10763,7.12589,7.14414,7.16239,7.18064,7.19889,7.21714,7.23539,7.25365,7.2719,7.29015,7.3084,7.32665,7.3449,7.36315,7.38141,7.39966,7.41791,7.43616,7.45441,7.47266,7.49091,7.50916,7.52742,7.54567,7.56392,7.58217,7.60042,7.61867,7.63692,7.65518,7.67343,7.69168,7.70993,7.72818,7.74643,7.76468,7.78293,7.80119,7.81944,7.83769,7.85594,7.87419,7.89244,7.91069,7.92895,7.9472,7.96545,7.9837,8.00195,8.0202,8.03845,8.05671,8.07496,8.09321,8.11146,8.12971,8.14796,8.16621,8.18446,8.20272,8.22097,8.23922,8.25747,8.27572,8.29397,8.31222,8.33048,8.34873,8.36698,8.38523,8.40348,8.42173,8.43998,8.45823,8.47649,8.49474,8.51299,8.53124,8.54949,8.56774,8.58599,8.60425,8.6225,8.64075,8.659,8.67725,8.6955,8.71375,8.732,8.75026,8.76851,8.78676,8.80501,8.82326,8.84151,8.85976,8.87802,8.89627,8.91452,8.93277,8.95102,8.96927,8.98752,9.00578,9.02403,9.04228,9.06053,9.07878,9.09703,9.11528,9.13353,9.15179,9.17004,9.18829,9.20654,9.22479,9.24304,9.26129,9.27955,9.2978,9.31605,9.3343,9.35255,9.3708,9.38905,9.4073,9.42556,9.44381,9.46206,9.48031,9.49856,9.51681,9.53506,9.55332,9.57157,9.58982,9.60807,9.62632,9.64457,9.66282,9.68108,9.69933,9.71758,9.73583,9.75408,9.77233,9.79058,9.80883,9.82709,9.84534,9.86359,9.88184,9.90009,9.91834,9.93659,9.95485,9.9731,9.99135,10.0096,10.0279,10.0461,10.0644,10.0826,10.1009,10.1191,10.1374,10.1556,10.1739,10.1921,10.2104,10.2286,10.2469,10.2651,10.2834,10.3016,10.3199,10.3381,10.3564,10.3746,10.3929,10.4111,10.4294,10.4476,10.4659,10.4841,10.5024,10.5206,10.5389,10.5571,10.5754,10.5936,10.6119,10.6301,10.6484,10.6666,10.6849,10.7032,10.7214,10.7397,10.7579,10.7762,10.7944,10.8127,10.8309,10.8492,10.8674,10.8857,10.9039,10.9222,10.9404,10.9587,10.9769,10.9952,11.0134,11.0317,11.0499,11.0682,11.0864,11.1047,11.1229,11.1412,11.1594,11.1777,11.1959,11.2142,11.2324,11.2507,11.2689,11.2872,11.3054,11.3237,11.3419,11.3602,11.3785,11.3967,11.415,11.4332,11.4515,11.4697,11.488,11.5062,11.5245,11.5427,11.561,11.5792,11.5975,11.6157,11.634,11.6522   ,11.6705,11.6887,11.707,11.7252,11.7435,11.7617,11.78,11.7982,11.8165,11.8347,11.853,11.8712,11.8895,11.9077,11.926,11.9442,11.9625,11.9807,11.999,12.0172,12.0355,12.0538,12.072,12.0903,12.1085,12.1268,12.145,12.1633,12.1815,12.1998,12.218,12.2363,12.2545,12.2728,12.291,12.3093,12.3275,12.3458,12.364,12.3823,12.4005,12.4188,12.437,12.4553,12.4735,12.4918,12.51,12.5283,12.5465,12.5648,12.583,12.6013,12.6195,12.6378,12.656,12.6743,12.6925,12.7108,12.7291,12.7473,12.7656,12.7838,12.8021,12.8203,12.8386,12.8568,12.8751,12.8933,12.9116,12.9298,12.9481,12.9663,12.9846,13.0028,13.0211,13.0393,13.0576,13.0758,13.0941,13.1123,13.1306,13.1488,13.1671,13.1853,13.2036,13.2218,13.2401,13.2583,13.2766,13.2948,13.3131,13.3313,13.3496,13.3678,13.3861,13.4044,13.4226,13.4409,13.4591,13.4774,13.4956,13.5139,13.5321,13.5504,13.5686,13.5869,13.6051,13.6234,13.6416,13.6599,13.6781,13.6964,13.7146,13.7329,13.7511,13.7694,13.7876,13.8059,13.8241,13.8424,13.8606,13.8789,13.8971,13.9154,13.9336,13.9519,13.9701,13.9884,14.0066,14.0249,14.0431,14.0614,14.0797,14.0979,14.1162,14.1344,14.1527,14.1709,14.1892,14.2074,14.2257,14.2439,14.2622,14.2804,14.2987,14.3169,14.3352,14.3534,14.3717,14.3899,14.4082,14.4264,14.4447,14.4629,14.4812,14.4994,14.5177,14.5359,14.5542,14.5724,14.5907,14.6089,14.6272,14.6454,14.6637,14.6819,14.7002,14.7184,14.7367,14.755,14.7732,14.7915,14.8097,14.828,14.8462,14.8645,14.8827,14.901,14.9192,14.9375,14.9557,14.974,14.9922,15.0105,15.047,15.0652,15.0835,15.12,15.1382,15.1565,15.1747,15.193,15.2112,15.2295,15.2477,15.266,15.2842,15.3025,15.3207,15.339,15.3572,15.3755,15.3937,15.412,15.4303,15.4485,15.4668,15.485,15.5033,15.5215,15.5398,15.558,15.5763,15.5945,15.6128,15.631,15.6493,15.6675,15.6858,15.704,15.7223,15.7405,15.7588,15.777,15.7953,15.8135,15.8318,15.85,15.8683,15.8865,15.9048,15.923,15.9413,15.9595,15.9778,15.996,16.0143,16.1421,16.1603,16.1786,16.1968,16.2151,16.2333,16.2516,16.2698,16.2881,16.3063,16.3246,16.3428,16.3611,16.3793,16.3976,16.4158,16.4341,16.4523,16.4706,16.4888,16.5071,16.5253,16.5436,16.5618,16.5801,16.5983,16.6166,16.6348,16.6531,16.6713,16.6896,16.7078,16.7261,16.7443,16.7626,16.7809,16.7991,16.8174,16.8356,16.8539,16.8721,16.8904,16.9086,16.9269,16.9451,16.9634,16.9816,16.9999,17.0181,17.0364,17.0546,17.0729,17.0911,17.1094,17.1276,17.1459,17.1641,17.1824,17.2006,17.2189,17.2371,17.2554,17.2736,17.2919,17.3101,17.3284,17.3466,17.3649,17.3831,17.4014,17.4196,17.4379,17.4562,17.4744,17.4927,17.5109,17.5292,17.5474,17.5657,17.5839,17.6022,17.6204,17.6387,17.6569,17.6752,17.6934,17.7117,17.7299,17.7482,17.7664,17.7847,17.8029,17.8212,17.8394,17.8577,17.8759,17.8942,17.9124,17.9307,17.9489,17.9672,17.9854,18.0037,18.0219,18.0402,18.0584,18.0767,18.0949,18.1132,18.1315,18.1497,18.168,18.1862,18.2045,18.2227,18.241,18.2592,18.2775,18.2957,18.314,18.3322,18.3505,18.3687,18.387,18.4052,18.4235,18.4417,18.46,18.4782,18.4965,18.5147,18.533,18.5512,18.5695,18.5877,18.606,18.6242,18.6425,18.6607,18.679,18.6972,18.7155,18.7337,18.752,18.7702,18.7885,18.8068,18.825,18.8433,18.8615,18.8798,18.898,18.9163,18.9345,18.9528,18.971,18.9893,19.0075,19.0258,19.044,19.0623,19.0805,19.0988,19.117,19.1353,19.1535,19.1718,19.19,19.2083,19.2265,19.2448,19.263,19.2813,19.2995,19.3178,19.336,19.3543,19.3725,19.3908,19.409,19.4273,19.4455,19.4638,19.4821,19.5003,19.5186,19.5368,19.5551,19.5733,19.5916,19.6098,19.6281,19.6463,19.6646,19.6828,19.7011,19.7193,19.7376,19.7558,19.7741,19.7923,19.8106,19.8288,19.8471,19.8653,19.8836,19.9018,19.9201,19.9383,19.9566,19.9748,19.9931,20.0113,20.0296,20.0478,20.0661,20.0843,20.1026,20.1208,20.1391,20.1574,20.1756,20.1939,20.2121,20.2304,20.2486,20.2669,20.2851,20.3034,20.3216,20.3399,20.3581,20.3764,20.3946,20.4129,20.4311,20.4494,20.4676,20.4859,20.5041,20.5224,20.5406,20.5589,20.5771,20.5954,20.6136,20.6319,20.6501,20.6684,20.6866,20.7049,20.7231,20.7414,20.7596,20.7779,20.7961,20.8144,20.8326,20.8509,20.8692,20.8874,20.9057,20.9239,20.9422,20.9604,20.9787,20.9969,21.0152,21.0334,21.0517,21.0699,21.0882,21.1064,21.1247,21.1429,21.1612,21.1794,21.1977,21.2159,21.2342,21.2524,21.2707,21.2889,21.3072,21.3254,21.3437,21.3619,21.3802,21.3984,21.4167,21.4349,21.4532,21.4714,21.4897,21.5079,21.5262,21.5445,21.5627,21.581,21.5992,21.6175,21.6357,21.654,21.6722,21.6905,21.7087,21.727,21.7452,21.7635,21.7817,21.8,21.8182,21.8365,21.8547,21.873,21.8912,21.9095,21.9277,21.946,21.9642,21.9825,22.0007,22.019,22.0372,22.0555,22.0737,22.092,22.1102,22.1285,22.1467,22.165,22.1832,22.2015,22.2198,22.238,22.2563,22.2745,22.2928,22.311,22.3293,22.3475,22.3658,22.384,22.4023,22.4205,22.4388,22.457,22.4753,22.4935,22.5118,22.53,22.5483,22.5665,22.5848,22.603,22.6213,22.6395,22.6578,22.676,22.6943,22.7125,22.7308,22.749,22.7673,22.7855,22.8038,22.822,22.8403,22.8585,22.8768,22.8951,22.9133,22.9316,22.9498,22.9681,22.9863,23.0046,23.0228,23.0411,23.0593,23.0776,23.0958,23.1141,23.1323,23.1506,23.1688,23.1871,23.2053,23.2236,23.2418,23.2601,23.2783,23.2966,23.3148,23.3331,23.3513,23.3696,23.3878,23.4061,23.4243,23.4426,23.4608,23.4791,23.4973,23.5156,23.5338,23.5521,23.5704,23.5886,23.6069,23.6251,23.6434,23.6616,23.6799,23.6981,23.7164,23.7346,23.7529,23.7711,23.7894,23.8076,23.8259,23.8441,23.8624,23.8806,23.8989,23.9171,23.9354,23.9536,23.9719,23.9901,24.0084,24.0266,24.0449,24.0631,24.0814,24.0996,24.1179,24.1361,24.1544,24.1726,24.1909,24.2091,24.2274,24.2457,24.2639,24.2822,24.3004,24.3187,24.3369,24.3552,24.3734,24.3917,24.4099,24.4282,24.4464,24.4647,24.4829,24.5012,24.5194,24.5377,24.5559,24.5742,24.5924,24.6107,24.6289,24.6472,24.6654,24.6837,24.7019,24.7202,24.7384,24.7567,24.7749,24.7932,24.8114,24.8297,24.8479,24.8662,24.8844,24.9027,24.921,24.9392,24.9575,24.9757,24.994,25.0122,25.0305,25.0487,25.067,25.0852,25.1035,25.1217,25.14,25.1582,25.1765,25.1947,25.213,25.2312,25.2495,25.2677,25.286,25.3042,25.3225,25.3407,25.359,25.3772,25.3955,25.4137,25.432,25.4502,25.4685,25.4867,25.505,25.5232,25.5415,25.5597,25.578,25.5963,25.6145,25.6328,25.651,25.6693,25.6875,25.7058,25.724,25.7423,25.7605,25.7788,25.797,25.8153,25.8335,25.8518,25.87,25.8883,25.9065,25.9248,25.943,25.9613,25.9795,25.9978,26.016,26.0343,26.0525,26.0708,26.089,26.1073,26.1255,26.1438,26.162,26.1803,26.1985,26.2168,26.235,26.2533,26.2716,26.2898,26.3081,26.3263,26.3446,26.3628,26.3811,26.3993,26.4176,26.4358,26.4541,26.4723,26.4906,26.5088,26.5271,26.5453,26.5636,26.5818,26.6001,26.6183,26.6366,26.6548,26.6731,26.6913,26.7096,26.7278,26.7461,26.7643,26.7826,26.8008,26.8191,26.8373,26.8556,26.8738,26.8921,26.9103,26.9286,26.9469,26.9651,26.9834,27.0016,27.0199,27.0381,27.0564,27.0746,27.0929,27.1111,27.1294,27.1476,27.1659,27.1841,27.2024,27.2206,27.2389,27.2571,27.2754,27.2936,27.3119,27.3301,27.3484,27.3666,27.3849,27.4031,27.4214,27.4396,27.4579,27.4761,27.4944,27.5126,27.5309,27.5491,27.5674,27.5856,27.6039,27.6222,27.6404,27.6587,27.6769,27.6952,27.7134,27.7317,27.7499,27.7682,27.7864,27.8047,27.8229,27.8412,27.8594,27.8777,27.8959,27.9142,27.9324,27.9507,27.9689,27.9872,28.0054,28.0237,28.0419,28.0602,28.0784,28.0967,28.1149,28.1332,28.1514,28.1697,28.1879,28.2062,28.2244,28.2427,28.2609,28.2792,28.2975,28.3157,28.334,28.3522,28.3705,28.3887,28.407,28.4252,28.4435,28.4617,28.48,28.4982,28.5165,28.5347,28.553,28.5712,28.5895,28.6077,28.626,28.6442,28.6625,28.6807,28.699,28.7172,28.7355,28.7537,28.772,28.7902,28.8085,28.8267,28.845,28.8632,28.8815,28.8997,28.918,28.9362,28.9545,28.9728,28.991,29.0093,29.0275,29.0458,29.064,29.0823,29.1005,29.1188,29.137,29.1553,29.1735,29.1918,29.21,29.2283,29.2465,29.2648,29.283,29.3013,29.3195,29.3378,29.356,29.3743,29.3925,29.4108,29.429,29.4473,29.4655,29.4838,29.502,29.5203,29.5385,29.5568,29.575,29.5933,29.6115,29.6298,29.6481,29.6663,29.6846,29.7028,29.7211,29.7393,29.7576,29.7758,29.7941,29.8123,29.8306,29.8488,29.8671,29.8853,29.9036,29.9218,29.9401,29.9583,29.9766,29.9948,30.0131,30.0313,30.0496,30.0678,30.0861,30.1043,30.1226,30.1408,30.1591,30.1773,30.1956,30.2138,30.2321,30.2503,30.2686,30.2868,30.3051,30.3234,30.3416,30.3599,30.3781,30.3964,30.4146,30.4329,30.4511,30.4694,30.4876,30.5059,30.5241,30.5424,30.5606,30.5789,30.5971,30.6154,30.6336,30.6519,30.6701,30.6884,30.7066,30.7249,30.7431,30.7614,30.7796,30.7979,30.8161,30.8344,30.8526,30.8709,30.8891,30.9074,30.9256,30.9439,30.9621,30.9804,30.9987,31.0169,31.0352,31.0534,31.0717,31.0899,31.1082,31.1264,31.1447,31.1629,31.1812,31.1994,31.2177,31.2359,31.2542,31.2724,31.2907,31.3089,31.3272,31.3454,31.3637,31.3819,31.4002,31.4184,31.4367,31.4549,31.4732,31.4914,31.5097,31.5279,31.5462,31.5644,31.5827,31.6009,31.6192,31.6374,31.6557,31.674,31.6922,31.7105,31.7287,31.747,31.7652,31.7835,31.8017,31.82,31.8382,31.8565,31.8747,31.893,31.9112,31.9295,31.9477,31.966,31.9842,32.0025,32.0207,32.039,32.0572,32.0755,32.0937,32.112,32.1302,32.1485,32.1667,32.185,32.2032,32.2215,32.2397,32.258,32.2762,32.2945,32.3127,32.331,32.3493,32.3675,32.3858,32.404,32.4223,32.4405,32.4588,32.477,32.4953,32.5135,32.5318,32.55,32.5683,32.5865,32.6048,32.623,32.6413,32.6595,32.6778,32.696,32.7143,32.7325,32.7508,32.769,32.7873,32.8055,32.8238,32.842,32.8603,32.8785,32.8968,32.915,32.9333,32.9515,32.9698,32.988,33.0063,33.0246,33.0428,33.0611,33.0793,33.0976,33.1158,33.1341,33.1523,33.1706,33.1888,33.2071,33.2253,33.2436,33.2618,33.2801,33.2983,33.3166,33.3348,33.3531,33.3713,33.3896,33.4078,33.4261,33.4443,33.4626,33.4808,33.4991,33.5173,33.5356,33.5538,33.5721,33.5903,33.6086,33.6268,33.6451,33.6633,33.6816,33.6999,33.7181,33.7364,33.7546,33.7729,33.7911,33.8094,33.8276,33.8459,33.8641,33.8824,33.9006,33.9189,33.9371,33.9554,33.9736,33.9919,34.0101,34.0284,34.0466,34.0649,34.0831,34.1014,34.1196,34.1379,34.1561,34.1744,34.1926,34.2109,34.2291,34.2474,34.2656,34.2839,34.3021,34.3204,34.3386,34.3569,34.3752,34.3934,34.4117,34.4299,34.4482,34.4664,34.4847,34.5029,34.5212,34.5394,34.5577,34.5759,34.5942,34.6124,34.6307,34.6489,34.6672,34.6854,34.7037,34.7219,34.7402,34.7584,34.7767,34.7949,34.8132,34.8314,34.8497,34.8679,34.8862,34.9044,34.9227,34.9409,34.9592,34.9774,34.9957,35.0139,35.0322,35.0505,35.0687,35.087,35.1052,35.1235,35.1417,35.16,35.1782,35.1965,35.2147,35.233,35.2512,35.2695,35.2877,35.306,35.3242,35.3425,35.3607,35.379,35.3972,35.4155,35.4337,35.452,35.4702,35.4885,35.5067,35.525,35.5432,35.5615,35.5797,35.598,35.6162,35.6345,35.6527,35.671,35.6892,35.7075,35.7258,35.744,35.7623,35.7805,35.7988,35.817,35.8353,35.8535,35.8718,35.89,35.9083,35.9265,35.9448,35.963,35.9813,35.9995,36.0178,36.036,36.0543,36.0725,36.0908,36.109,36.1273,36.1455,36.1638,36.182,36.2003,36.2185,36.2368,36.255,36.2733,36.2915,36.3098,36.328,36.3463,36.3645,36.3828,36.4011,36.4193,36.4376,36.4558,36.4741,36.4923,36.5106,36.5288,36.5471,36.5653,36.5836,36.6018,36.6201,36.6383,36.6566,36.6748,36.6931,36.7113,36.7296,36.7478,36.7661,36.7843,36.8026,36.8208,36.8391,36.8573,36.8756,36.8938,36.9121,36.9303,36.9486,36.9668,36.9851,37.0033,37.0216,37.0398,37.0581,37.0764,37.0946,37.1129,37.1311,37.1494,37.1676,37.1859,37.2041,37.2224,37.2406,37.2589,37.2771,37.2954,37.3136,37.3319,37.3501,37.3684,37.3866,37.4049,37.4231,37.4414,37.4596,37.4779,37.4961,37.5144,37.5326,37.5509,37.5691,37.5874,37.6056,37.6239,37.6421,37.6604,37.6786,37.6969,37.7151,37.7334,37.7517,37.7699,37.7882,37.8064,37.8247,37.8429,37.8612,37.8794,37.8977,37.9159,37.9342,37.9524,37.9707,37.9889,38.0072,38.0254,38.0437,38.0619,38.0802,38.0984,38.1167,38.1349,38.1532,38.1714,38.1897,38.2079,38.2262,38.2444,38.2627,38.2809,38.2992,38.3174,38.3357,38.3539,38.3722,38.3904,38.4087,38.427,38.4452,38.4635,38.4817,38.5,38.5182,38.5365,38.5547,38.573,38.5912,38.6095,38.6277,38.646,38.6642,38.6825,38.7007,38.719,38.7372,38.7555,38.7737,38.792,38.8102,38.8285,38.8467,38.865,38.8832,38.9015,38.9197,38.938,38.9562,38.9745,38.9927,39.011,39.0292,39.0475,39.0657,39.084;

idx_rfr_saharan_dust_rl = 1.53,
1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,1.56,
1.560000,1.559800,1.559900,1.559800,1.551800,1.550100,
1.4529,1.45264,1.45237,1.45207,1.45626,1.45554,1.45918,1.45947,1.45896,1.4623,1.46321,1.46707,1.46656,1.4663,1.46584,1.4685,1.46974,1.46815,1.46764,1.46487,1.46447,1.46428,1.46401,1.46375,1.46324,1.4669,1.46781,1.47113,1.47373,1.4789,1.48111,1.48696,1.49003,1.4951,1.50041,1.50264,1.5022,1.50193,1.50167,1.50144,1.49531,1.49293,1.48329,1.47715,1.4754,1.46632,1.46075,1.4576,1.45715,1.45972,1.46106,1.4606,1.4628,1.46453,1.46416,1.46395,1.46374,1.46338,1.46505,1.4671,1.47102,1.47076,1.47057,1.4703,1.47004,1.46977,1.46946,1.47366,1.47294,1.47675,1.47317,1.47685,1.47634,1.47607,1.47581,1.47554,1.47522,1.47676,1.47913,1.47878,1.48287,1.48237,1.48211,1.48179,1.48405,1.4856,1.48537,1.48486,1.48821,1.48878,1.48851,1.48825,1.48798,1.48772,1.48745,1.48719,1.48692,1.48666,1.4864,1.48624,1.48596,1.4857,1.48525,1.48781,1.48916,1.48977,1.49303,1.49225,1.50076,1.50031,1.49991,1.50401,1.50373,1.5033,1.50718,1.50715,1.5067,1.51032,1.51056,1.51035,1.51014,1.51038,1.514,1.51355,1.51352,1.5172,1.51968,1.52078,1.52481,1.52676,1.52837,1.53293,1.53617,1.54167,1.54406,1.55238,1.5559,1.55994,1.56808,1.5741,1.58222,1.59016,1.5963,1.60056,1.60009,1.60011,1.58901,1.56809,1.55453,1.54222,1.52777,1.50799,1.49571,1.48926,1.48046,1.47441,1.46841,1.46313,1.45835,1.45405,1.45308,1.44962,1.4453,1.44503,1.44198,1.44023,1.43545,1.43547,1.43521,1.43514,1.43198,1.43029,1.43004,1.42977,1.42951,1.42925,1.42898,1.42862,1.43299,1.43012,1.42783,1.43214,1.4317,1.43144,1.43061,1.42641,1.42627,1.4305,1.43037,1.42655,1.42548,1.42521,1.42495,1.42468,1.42467,1.42094,1.41978,1.41952,1.41925,1.41899,1.41872,1.41846,1.41819,1.41796,1.41777,1.4175,1.41724,1.41697,1.4167,1.41644,1.41618,1.41591,1.41564,1.41544,1.41522,1.41495,1.41469,1.41442,1.41416,1.41389,1.41363,1.41336,1.41315,1.41294,1.41315,1.4168,1.41636,1.41605,1.41733,1.41996,1.4195,1.42042,1.42316,1.42656,1.42678,1.42636,1.42951,1.43447,1.4339,1.43683,1.4378,1.43878,1.44145,1.44501,1.44592,1.44935,1.44866,1.45288,1.45252,1.45225,1.45199,1.45172,1.45146,1.4512,1.45093,1.45073,1.45052,1.44734,1.44731,1.4455,1.4393,1.43647,1.43589,1.42746,1.42416,1.41807,1.41197,1.40599,1.39995,1.39419,1.38411,1.37971,1.37142,1.36421,1.35125,1.34861,1.33862,1.32821,1.32032,1.31529,1.30477,1.29506,1.28935,1.27672,1.26835,1.26168,1.24882,1.24176,1.23324,1.22917,1.21764,1.20862,1.20232,1.19461,1.18663,1.18376,1.17407,1.16845,1.16682,1.16056,1.15451,1.14852,1.14243,1.13645,1.13036,1.12438,1.1181,1.11617,1.106,1.09999,1.09844,1.08912,1.09005,1.08069,1.07905,1.07261,1.07188,1.06969,1.06331,1.06184,1.05821,1.05397,1.05355,1.05358,1.04902,1.04839,1.05068,1.05231,1.05174,1.05511,1.06559,1.07536,1.09329,1.11348,1.14597,1.17689,1.22532,1.30264,1.38057,1.42693,1.45127,1.49094,1.55463,1.54141,1.59183,1.70822,1.76198,1.77635,1.81618,1.83904,1.84817,1.85324,1.8596,1.87458,1.89342,1.91532,1.93429,1.95349,1.99517,2.07046,2.13625,2.16891,2.2063,2.23525,2.30465,2.37685,2.43263,2.48099,2.527,2.57085,2.61661,2.66245,2.70069,2.74143,2.77705,2.80653,2.84703,2.88426,2.90868,2.92736,2.95346,2.97869,2.99297,3.00569,3.01564,3.02178,3.02604,3.02594,3.02173,3.01456,3.00178,2.99397,2.97041,2.95516,2.93153,2.91683,2.88861,2.86172,2.82834,2.79689,2.76196,2.73776,2.70735,2.68009,2.65252,2.61922,2.5926,2.56153,2.5302,2.5061,2.47724,2.45778,2.42248,2.39074,2.36638,2.33483,2.29458,2.25206,2.21814,2.17314,2.13909,2.10185,2.07171,2.04827,2.03271,2.00855,1.98192,1.94813,1.92771,1.88735,1.8504,1.81442,1.78302,1.77478,1.75021,1.73177,1.71934,1.71271,1.70681,1.70068,1.69914,1.69562,1.69561,1.69617,1.70347,1.71385,1.71987,1.73057,1.7436,1.75324,1.76318,1.77306,1.78301,1.79316,1.80032,1.80547,1.81367,1.81271,1.81637,1.821,1.82061,1.82016,1.82444,1.82839,1.82787,1.8277,1.82744,1.82788,1.81827,1.81833,1.81807,1.81784,1.81303,1.81327,1.80865,1.80842,1.80816,1.8079,1.80763,1.80736,1.8071,1.80687,1.80667,1.8064,1.80614,1.80588,1.80561,1.80535,1.80509,1.80483,1.80361,1.79997,1.79991,1.79965,1.79969,1.79538,1.79475,1.79448,1.79422,1.79409,1.79127,1.78917,1.78906,1.78879,1.78871,1.78381,1.78378,1.78352,1.78328,1.7831,1.78282,1.78256,1.7826,1.77834,1.77758,1.7774,1.77713,1.7762,1.7721,1.77213,1.77196,1.76947,1.76715,1.76711,1.76441,1.76222,1.76206,1.7618,1.76171,1.7568,1.75709,1.75276,1.75216,1.7519,1.75162,1.75054,1.74671,1.74672,1.74571,1.7417,1.74173,1.74056,1.73687,1.73682,1.73656,1.7363,1.73602,1.73576,1.73549,1.73532,1.73506,1.73454,1.73813,1.73417,1.73401,1.73375,1.73376,1.73769,1.73716,1.73689,1.73662,1.73643,1.73621,1.73593,1.73567,1.73541,1.73515,1.73487,1.73461,1.73435,1.73408,1.73403,1.72916,1.72949,1.72482,1.72475,1.72163,1.71984,1.71507,1.71548,1.71069,1.70889,1.70896,1.70567,1.70715,1.70685,1.70498,1.70473,1.70447,1.70421,1.70394,1.70367,1.70351,1.70325,1.70298,1.70272,1.70246,1.7025,1.69812,1.6967,1.69281,1.69281,1.69146,1.68823,1.68369,1.68366,1.68065,1.6745,1.67433,1.67436,1.66946,1.66491,1.66523,1.66052,1.65852,1.65568,1.65513,1.64891,1.64661,1.64581,1.6395,1.63754,1.63754,1.63473,1.62868,1.62846,1.62513,1.62351,1.61883,1.61887,1.6186,1.61734,1.61077,1.60952,1.60776,1.6049,1.60027,1.60033,1.59682,1.5911,1.59101,1.59074,1.59009,1.58361,1.58152,1.58137,1.58139,1.57733,1.57657,1.57395,1.57166,1.57059,1.56712,1.56277,1.56235,1.56209,1.56182,1.5607,1.55697,1.55702,1.55218,1.55228,1.55215,1.54727,1.5475,1.54304,1.54263,1.54237,1.5422,1.53757,1.53457,1.533,1.53292,1.52957,1.52781,1.52339,1.52389,1.5145,1.51451,1.51471,1.50379,1.48724,1.48884,1.50575,1.51041,1.51373,1.50917,1.49868,1.49776,1.49687,1.49603,1.49526,1.49459,1.49431,1.49441,1.49454,1.49461,1.49456,1.49431,1.49312,1.49149,1.48976,1.48804,1.48644,1.48542,1.48519,1.48515,1.48522,1.48533,1.4854,1.48501,1.48434,1.48358,1.48275,1.48187,1.48097,1.48007,1.47918,1.47835,1.47759,1.47693,1.47654,1.47638,1.47631,1.47633,1.47639,1.47648,1.47672,1.47693,1.47706,1.47703,1.47681,1.47626,1.47475,1.47307,1.46718,1.46738,1.4676,1.46758,1.46756,1.46755,1.46753,1.46751,1.46749,1.46746,1.46743,1.46739,1.46735,1.46732,1.46721,1.46708,1.46698,1.46693,1.46695,1.46707,1.46759,1.46826,1.46898,1.46971,1.4704,1.47102,1.47113,1.47109,1.471,1.47092,1.47087,1.47093,1.47133,1.47184,1.47246,1.47321,1.47406,1.47506,1.47634,1.47769,1.47908,1.48046,1.48181,1.48309,1.48345,1.4838,1.48426,1.48491,1.48587,1.48726,1.49074,1.49472,1.49909,1.50373,1.50854,1.51341,1.51822,1.52196,1.52473,1.52747,1.53028,1.53326,1.5365,1.54011,1.54582,1.55274,1.56016,1.56796,1.57605,1.58432,1.59265,1.60095,1.6091,1.617,1.62454,1.63161,1.63811,1.64394,1.64897,1.65312,1.65626,1.65953,1.67091,1.68322,1.69635,1.71016,1.72455,1.73939,1.75456,1.76995,1.78543,1.80089,1.8162,1.83125,1.84592,1.86008,1.87363,1.88643,1.89837,1.90933,1.9192,1.92296,1.92533,1.92826,1.93172,1.93567,1.94008,1.94491,1.95013,1.95571,1.9616,1.96777,1.97419,1.98083,1.98764,1.9946,2.0017,2.00916,2.01663,2.02405,2.03137,2.03851,2.04542,2.05204,2.05831,2.0637,2.06581,2.06798,2.07045,2.07352,2.07743,2.08246,2.08948,2.10664,2.1256,2.14584,2.16686,2.18817,2.20925,2.22961,2.24874,2.26614,2.27899,2.28481,2.28902,2.2918,2.29336,2.29388,2.29355,2.29294,2.29193,2.29043,2.28853,2.28631,2.28404,2.28185,2.27949,2.27694,2.27421,2.27118,2.26773,2.26418,2.26062,2.25713,2.25405,2.25153,2.2491,2.24669,2.24421,2.24135,2.23779,2.2342,2.23066,2.2273,2.22456,2.22259,2.2209,2.2194,2.21805,2.21669,2.21486,2.21308,2.21142,2.20992,2.20863,2.20812,2.20797,2.20798,2.20807,2.20817,2.20816,2.20732,2.20642,2.20553,2.20471,2.20405,2.20387,2.20419,2.20474,2.20548,2.20639,2.20744,2.20857,2.20976,2.21103,2.21237,2.21374,2.21515,2.21646,2.2176,2.2188,2.22006,2.22142,2.22291,2.22469,2.2271,2.22963,2.23223,2.23483,2.23738,2.23982,2.24165,2.24301,2.24429,2.24554,2.24682,2.24818,2.24991,2.25208,2.25442,2.2569,2.25952,2.26224,2.26507,2.26794,2.27087,2.27386,2.2769,2.27997,2.28307,2.28619,2.28894,2.29173,2.2946,2.29759,2.30075,2.30412,2.30789,2.31264,2.31765,2.32286,2.32821,2.33366,2.33914,2.34462,2.34985,2.35444,2.35895,2.36341,2.36784,2.37225,2.37666,2.3811,2.38577,2.39055,2.39537,2.40022,2.4051,2.41,2.41492,2.41985,2.4248,2.42976,2.43469,2.43961,2.4445,2.44935,2.45415,2.45884,2.46337,2.46786,2.47231,2.47672,2.48111,2.48548,2.48985,2.49441,2.49898,2.50352,2.50802,2.51245,2.51681,2.52106,2.52501,2.52851,2.53197,2.53542,2.53891,2.54249,2.54621,2.55037,2.55523,2.56028,2.56549,2.5708,2.5762,2.58164,2.58709,2.59219,2.5968,2.60143,2.60612,2.61092,2.61586,2.62099,2.62635,2.63299,2.64027,2.64778,2.65545,2.66321,2.671,2.67875,2.68638,2.69383,2.70082,2.70707,2.71302,2.71867,2.72401,2.72902,2.73368,2.73798,2.74158,2.74432,2.74684,2.74924,2.7516,2.75401,2.75655,2.7599,2.76367,2.76771,2.77202,2.7766,2.78146,2.78659,2.79216,2.79844,2.80495,2.81162,2.81841,2.82527,2.83213,2.83894,2.84565,2.85178,2.85736,2.86281,2.86812,2.87333,2.87843,2.88346,2.88842,2.89358,2.89886,2.90405,2.90911,2.91403,2.91877,2.92331,2.92761,2.93109,2.9343,2.93736,2.94031,2.9432,2.94607,2.949,2.95241,2.95589,2.95943,2.963,2.96661,2.97023,2.97386,2.97749,2.9811,2.98469,2.98825,2.99177,2.99523,2.99862,3.00178,3.00486,3.0079,3.0109,3.01387,3.01683,3.0198,3.02295,3.02609,3.0292,3.03228,3.03531,3.03827,3.04116,3.04396,3.04666,3.04924,3.05168,3.05398,3.05611,3.05802,3.05973,3.06124,3.06255,3.06366,3.06455,3.06508,3.06528,3.06533,3.06524,3.06508,3.06486,3.06478,3.06474,3.06471,3.06467,3.06464,3.0646,3.06457,3.06453,3.0645,3.06446,3.06443,3.06446,3.06469,3.06485,3.06489,3.06477,3.06443,3.06354,3.06218,3.06061,3.0589,3.0571,3.05535,3.05387,3.05236,3.05077,3.04907,3.04724,3.04485,3.04233,3.03977,3.03724,3.0348,3.033,3.03142,3.02989,3.02835,3.02673,3.02473,3.02235,3.01985,3.01727,3.01464,3.0122,3.01003,3.00774,3.00526,3.00248,2.99905,2.9947,2.99011,2.98544,2.98081,2.97679,2.97319,2.96974,2.96638,2.96308,2.95942,2.95571,2.95212,2.94875,2.94565,2.94376,2.94221,2.94077,2.9393,2.93764,2.9351,2.93187,2.9284,2.92476,2.92103,2.91739,2.91382,2.91031,2.90691,2.90365,2.90082,2.89822,2.89574,2.89335,2.891,2.88868,2.88632,2.8839,2.88138,2.87871,2.87558,2.87211,2.86857,2.86505,2.86162,2.85868,2.85605,2.85354,2.85112,2.84877,2.84624,2.84362,2.84107,2.8386,2.83624,2.83448,2.83319,2.83185,2.83031,2.82841,2.82571,2.82138,2.81676,2.81205,2.80743,2.80375,2.80093,2.79841,2.79611,2.79393,2.79164,2.78915,2.78666,2.78416,2.78167,2.77917,2.77665,2.77414,2.77163,2.76912,2.76661,2.76411,2.76162,2.75913,2.75664,2.75412,2.7515,2.74891,2.7464,2.74399,2.74176,2.74025,2.7388,2.73731,2.73567,2.73378,2.73067,2.72707,2.72344,2.71993,2.71672,2.71527,2.71438,2.71373,2.71317,2.71253,2.71117,2.70873,2.70614,2.70353,2.70101,2.69902,2.69812,2.69741,2.69676,2.69604,2.69513,2.69339,2.69121,2.68876,2.68606,2.68314,2.67981,2.67626,2.67271,2.66927,2.66603,2.66379,2.66204,2.66047,2.65899,2.65749,2.65557,2.65321,2.65074,2.64818,2.64557,2.64294,2.64032,2.63775,2.63525,2.63287,2.63076,2.62911,2.62754,2.62599,2.62441,2.62271,2.62029,2.61777,2.61521,2.61268,2.61024,2.60847,2.60687,2.60533,2.60377,2.60212,2.6 ,2.59751,2.59496,2.59241,2.58992,2.58785,2.58622,2.58466,2.58311,2.58151,2.57967,2.57711,2.57449,2.57191,2.56946,2.5673,2.56621,2.56536,2.56465,2.56401,2.56334,2.56233,2.56099,2.5595,2.55784,2.55602,2.55396,2.55151,2.54897,2.54641,2.5439,2.54154,2.53972,2.53803,2.53645,2.53494,2.53346,2.53178,2.53008,2.52842,2.52685,2.52538,2.52425,2.52343,2.52269,2.52196,2.52119,2.52033,2.51894,2.51742,2.5158,2.51412,2.5124,2.51074,2.50912,2.5075,2.50588,2.50426,2.50265,2.50105,2.49945,2.49786,2.49626,2.49466,2.49304,2.49142,2.4898,2.48818,2.48656,2.48496,2.48336,2.48176,2.48016,2.47856,2.47696,2.47534,2.47372,2.4721,2.47048,2.46885,2.46701,2.46523,2.46356,2.46206,2.46076,2.46034,2.46031,2.4604,2.46049,2.46049,2.46028,2.45902,2.45753,2.45588,2.4541,2.45226,2.45041,2.4486,2.44688,2.44531,2.44393,2.44304,2.44281,2.44276,2.44283,2.44293,2.443,2.4426,2.44193,2.44117,2.44034,2.43946,2.43858,2.43779,2.43699,2.4362,2.4354,2.4346,2.43381,2.43301,2.43221,2.43142,2.43062,2.42983,2.42905,2.42828,2.4275,2.42673,2.42595,2.42516,2.42437,2.42358,2.42278,2.42198,2.42118,2.42027,2.41938,2.41853,2.41777,2.4171,2.41674,2.4167,2.41673,2.41678,2.4168,2.41674,2.41627,2.41558,2.41479,2.41394,2.41304,2.41212,2.4112,2.41032,2.40949,2.40874,2.40809,2.40774,2.40761,2.40757,2.4076,2.40768,2.40779,2.40802,2.40821,2.40831,2.40825,2.40798,2.4073,2.40576,2.40407,2.40234,2.40066,2.39914,2.39859,2.39837,2.39834,2.39847,2.39868,2.3989,2.39886,2.39883,2.3988,2.39876,2.39872,2.39869,2.39865,2.39862,2.39858,2.39855,2.39851,2.39848,2.39844,2.3984,2.39837,2.39833,2.3983,2.39828,2.39827,2.39825,2.39823,2.39822,2.3982,2.39817,2.39813,2.3981,2.39806,2.39802,2.39799,2.39795,2.39792,2.39788,2.39785,2.39781,2.39778,2.39774,2.3977,2.39767,2.39763,2.3976,2.39758,2.39757,2.39755,2.39753,2.39752,2.39749,2.39746,2.39743,2.3974,2.39736,2.39732,2.39729,2.39725,2.39722,2.39718,2.39715,2.39711,2.39707,2.39704,2.397,2.39697,2.39693,2.3969,2.39688,2.39687,2.39685,2.39683,2.39682,2.39678,2.39664,2.39652,2.39644,2.39643,2.39651,2.39684,2.39748,2.39818,2.39891,2.39962,2.40028,2.40062,2.40061,2.40054,2.40045,2.40038,2.40038,2.40083,2.4015,2.40221,2.40294,2.40364,2.40427,2.40453,2.4046,2.4046,2.40453,2.40443,2.4043,2.40427,2.40424,2.4042,2.40416,2.40413,2.40406,2.40392,2.4038,2.40373,2.40373,2.40382,2.40419,2.40484,2.40555,2.40628,2.40699,2.40763,2.40792,2.4079,2.40783,2.40774,2.40768,2.40768,2.40817,2.40884,2.40956,2.4103,2.411,2.41162,2.41184,2.41191,2.4119,2.41183,2.41172,2.41158,2.41144,2.41132,2.41125,2.41123,2.4113,2.41161,2.41224,2.41294,2.41367,2.41439,2.41504,2.41547,2.41556,2.41556,2.4155,2.41539,2.41525,2.41519,2.41517,2.41515,2.41514,2.41512,2.4151,2.41497,2.41485,2.41476,2.41473,2.41477,2.41497,2.41559,2.41629,2.41703,2.41775,2.41843,2.41894,2.41906,2.41908,2.41902,2.41892,2.41878,2.41868,2.41865,2.41861,2.41857,2.41854,2.41851,2.41841,2.41829,2.41821,2.41819,2.41824,2.41839,2.41898,2.41966,2.42038,2.42111,2.42179,2.42239,2.42254,2.42258,2.42254,2.42244,2.42231,2.42219,2.42216,2.42212,2.42209,2.42205,2.42202,2.42198,2.42194,2.42191,2.42187,2.42184,2.42181,2.42188,2.42197,2.42203,2.42201,2.42191,2.42168,2.42096,2.42014,2.41929,2.41845,2.41766,2.41717,2.41699,2.41692,2.41692,2.41698,2.41707,2.41709,2.41707,2.41705,2.41704,2.41702,2.417,2.41697,2.41694,2.4169,2.41687,2.41683,2.41679,2.41676,2.41672,2.41669,2.41665,2.41662,2.41658,2.41655,2.41651,2.41648,2.41644,2.41641,2.41647,2.41654,2.41658,2.41655,2.41644,2.41621,2.4155,2.41469,2.41385,2.41302,2.41225,2.41177,2.4116,2.41153,2.41153,2.41159,2.41168,2.41167,2.41163,2.4116,2.41156,2.41153,2.4115,2.41161,2.41169,2.41173,2.4117,2.41158,2.41124,2.41049,2.40966,2.40881,2.40797,2.40721,2.40682,2.40667,2.40662,2.40664,2.4067,2.40679,2.40676,2.40673,2.40669,2.40666,2.40662,2.4066,2.40658,2.40656,2.40654,2.40653,2.40651,2.40649,2.40646,2.40642,2.40639,2.40635,2.40631,2.40636,2.40644,2.40647,2.40644,2.40633,2.4061,2.40539,2.4046,2.40377,2.40294,2.40218,2.40168,2.40151,2.40143,2.40143,2.40149,2.40157,2.40167,2.40174,2.40178,2.40176,2.40164,2.40141,2.4007,2.39989,2.39904,2.3982,2.39741,2.39689,2.39673,2.39667,2.39669,2.39676,2.39686,2.39688,2.39685,2.39681,2.39678,2.39674,2.3967,2.39667,2.39663,2.3966,2.39656,2.39653,2.39651,2.3966,2.39667,2.39668,2.39661,2.39645,2.39602,2.39526,2.39443,2.39359,2.39278,2.39205,2.39178,2.39166,2.39162,2.39165,2.39172,2.39182,2.3919,2.39196,2.39197,2.39191,2.39175,2.39131,2.39056,2.38974,2.38891,2.3881,2.38738,2.38709,2.38696,2.38692,2.38695,2.38702,2.3871,2.38706,2.38703,2.38699,2.38696,2.38692,2.38694,2.38702,2.38707,2.38707,2.38698,2.3868,2.38634,2.38568,2.38492,2.38409,2.38322,2.38232,2.38141,2.38052,2.37968,2.37892,2.37826,2.37785,2.37769,2.37762,2.37763,2.37769,2.37779,2.37802,2.37823,2.37835,2.37833,2.37811,2.37755,2.37604,2.37436,2.37262,2.37093,2.36939,2.36871,2.36845,2.36838,2.36847,2.36867,2.3689,2.36901,2.3691,2.36913,2.3691,2.36897,2.3686,2.36785,2.36702,2.36616,2.36533,2.36457,2.36393,2.36346,2.3632,2.36321,2.36352,2.3642  ;

idx_rfr_saharan_dust_img = 0.070,
0.050561,0.045743,0.038785,0.031728,0.027208,0.023094,0.019765,0.016975,0.014397,0.012447,0.010859,0.009481,0.008340,0.007342,0.006425,0.005638,0.004929,0.004435,0.003992,0.003811,0.003810,0.003774,0.003773,
0.003300,0.003400,0.003600,0.003900,0.005600,0.005100,
0.017013,0.018438,0.019129,0.022541,0.027046,0.027542,0.027738,0.029433,0.032607,0.034432,0.034717,0.034863,0.034814,0.034415,0.034118,0.033743,0.033044,0.032163,0.029886,0.026572,0.023714,0.022342,0.022895,0.029880,0.021655,0.016871,0.016988,0.016101,0.015513,0.014854,0.014766,0.014771,0.014618,0.014386,0.014275,0.014029,0.013873,0.013794,0.013616,0.013436,0.013409,0.013316,0.013240,0.013096,0.012844,0.012617,0.012276,0.012017,0.011884,0.011805,0.011739,0.011608,0.011451,0.011160,0.010982,0.010837,0.010608,0.010430,0.010193,0.009949,0.009524,0.009204,0.008906,0.008288,0.008259,0.006893,0.006256,0.004783,0.004980,0.005012,0.004471,0.004473,0.004363,0.004307,0.004309,0.004286,0.004266,0.004305,0.004276,0.004286,0.004292,0.004302,0.004307,0.004353,0.004397,0.004443,0.004489,0.004533,0.004602,0.004669,0.004716,0.004774,0.004948,0.005082,0.005083,0.005270,0.005527,0.005679,0.005762,0.005817,0.005932,0.006055,0.006177,0.006333,0.006691,0.006928,0.007300,0.007507,0.007690,0.007759,0.007936,0.008439,0.008894,0.009233,0.009910,0.010280,0.010576,0.010876,0.011198,0.011673,0.012185,0.013203,0.013453,0.013654,0.013894,0.014060,0.014352,0.014641,0.015030,0.015506,0.015836,0.016224,0.016995,0.017693,0.017935,0.018441,0.018607,0.018989,0.019333,0.019691,0.020120,0.020762,0.021289,0.021843,0.023114,0.023852,0.024423,0.024928,0.025361,0.025618,0.026096,0.026440,0.027160,0.028022,0.028636,0.029519,0.030561,0.031870,0.032667,0.033312,0.033631,0.034173,0.034394,0.034990,0.035713,0.036451,0.037205,0.037973,0.038714,0.039049,0.040462,0.040711,0.041353,0.042553,0.042966,0.043432,0.043547,0.043937,0.044305,0.044254,0.044529,0.044998,0.045798,0.046084,0.046572,0.046858,0.047764,0.048611,0.049900,0.049745,0.050592,0.050617,0.050792,0.051066,0.051051,0.050581,0.050608,0.050407,0.049050,0.048795,0.047173,0.046188,0.045018,0.044007,0.043066,0.042106,0.041865,0.041876,0.042710,0.045052,0.046888,0.047116,0.048958,0.051981,0.056055,0.061754,0.066753,0.069496,0.071746,0.071110,0.057902,0.094201,0.086592,0.088522,0.092026,0.094634,0.100149,0.102806,0.103776,0.104558,0.104971,0.106149,0.10629,0.106267,0.106307,0.105574,0.105314,0.105199,0.103678,0.101258,0.101659,0.100856,0.100148,0.099129,0.097617,0.095271,0.091714,0.090449,0.088781,0.086347,0.085810,0.084481,0.082192,0.080417,0.078370,0.076275,0.075358,0.072422,0.071028,0.068546,0.066224,0.065525,0.064791,0.064560,0.063990,0.063411,0.063429,0.063418,0.063407,0.063470,0.064176,0.064457,0.064910,0.065591,0.066242,0.067249,0.068232,0.068907,0.070235,0.070899,0.072051,0.073028,0.073793,0.075334,0.076890,0.078561,0.078823,0.081817,0.083181,0.084928,0.085804,0.087266,0.089185,0.092035,0.094448,0.095584,0.098292,0.100674,0.10509,0.1076,0.108568,0.110659,0.114265,0.122015,0.125828,0.131309,0.135701,0.13929,0.141691,0.146168,0.151962,0.155577,0.163761,0.171838,0.175816,0.177372,0.180874,0.185595,0.191849,0.195619,0.199675,0.205241,0.222609,0.233777,0.244524,0.252867,0.253985,0.264424,0.277892,0.306018,0.320842,0.326846,0.337086,0.346595,0.351276,0.360086,0.371105,0.376641,0.396459,0.412026,0.423363,0.428527,0.432777,0.439112,0.448633,0.454073,0.459236,0.46889,0.478584,0.488491,0.498568,0.509078,0.517714,0.522484,0.532361,0.533428,0.538829,0.547573,0.551012,0.560564,0.561352,0.567685,0.5695,0.578564,0.589515,0.592256,0.605154,0.617649,0.630448,0.636939,0.64347,0.649762,0.661997,0.664067,0.674279,0.679787,0.695166,0.697174,0.710568,0.717247,0.729089,0.737945,0.772807,0.784678,0.791219,0.797860,0.804065,0.813336,0.831251,0.839201,0.844646,0.853808,0.871996,0.886437,0.894222,0.918693,0.929136,0.939144,0.943991,0.943391,0.942237,0.92733,0.913961,0.896719,0.887175,0.868527,0.845313,0.824644,0.80013,0.789922,0.772608,0.7567,0.740758,0.733402,0.721708,0.705693,0.691852,0.680581,0.661703,0.6477,0.633351,0.600296,0.5757,0.5642,0.552278,0.542367,0.53701,0.526689,0.519232,0.508355,0.502544,0.491719,0.481946,0.475394,0.465349,0.447007,0.440962,0.426193,0.41821,0.413736,0.406762,0.405737,0.395369,0.392975,0.384495,0.379883,0.375216,0.366727,0.36101,0.354893,0.343715,0.339451,0.329435,0.322122,0.320028,0.314479,0.313046,0.309062,0.304971,0.303606,0.297802,0.294736,0.291565,0.288535,0.28249,0.273923,0.26543,0.264521,0.257195,0.254617,0.252103,0.2471,0.247215,0.246222,0.243504,0.238833,0.233619,0.228668,0.223611,0.222896,0.218989,0.217258,0.215354,0.211702,0.211307,0.208915,0.206749,0.204446,0.203813,0.200052,0.197786,0.199024,0.197182,0.194922,0.193936,0.193982,0.193956,0.19375,0.195889,0.195949,0.195478,0.195441,0.19541,0.195377,0.19534,0.195221,0.190544,0.187003,0.183924,0.1807,0.180134,0.178186,0.174872,0.171619,0.170314,0.168583,0.168692,0.168249,0.165744,0.163901,0.162963,0.160134,0.159158,0.156457,0.154955,0.15197,0.15214,0.151291,0.149654,0.146873,0.146062,0.14359,0.142082,0.14057,0.13946,0.138755,0.138206,0.1382,0.136945,0.136851,0.138672,0.140443,0.141836,0.143788,0.146102,0.147522,0.149029,0.148842,0.150148,0.153562,0.154028,0.156965,0.158434,0.160989,0.163133,0.166257,0.167807,0.171066,0.174456,0.176041,0.181461,0.186145,0.187854,0.189781,0.191716,0.193703,0.195783,0.19768,0.201447,0.201534,0.202078,0.204366,0.204895,0.206831,0.208487,0.208232,0.209549,0.211796,0.211814,0.211776,0.21174,0.211829,0.207919,0.208277,0.205705,0.20441,0.204447,0.204505,0.203461,0.201119,0.200859,0.200821,0.201001,0.198124,0.197339,0.197302,0.197381,0.195976,0.195523,0.195443,0.19613,0.197189,0.197105,0.19531,0.19533,0.195291,0.195196,0.196928,0.19679,0.197544,0.19985,0.200143,0.200047,0.200683,0.202966,0.203453,0.203357,0.20388,0.206187,0.206843,0.206961,0.210414,0.210225,0.210188,0.21012,0.211939,0.212661,0.213741,0.213614,0.213577,0.213539,0.213502,0.213466,0.213429,0.213391,0.213354,0.213216,0.21505,0.215074,0.214928,0.216375,0.21516,0.215215,0.216835,0.216682,0.216645,0.216609,0.21657,0.216534,0.216399,0.218278,0.218198,0.219127,0.220155,0.220033,0.219995,0.219947,0.219911,0.219875,0.219836,0.2198,0.219763,0.219727,0.219707,0.219159,0.217771,0.216284,0.215839,0.215741,0.216557,0.217546,0.21924,0.221253,0.221857,0.223151,0.223006,0.222967,0.22292,0.222885,0.222846,0.22281,0.222704,0.223296,0.222643,0.222574,0.224557,0.224346,0.226341,0.226067,0.22829,0.230197,0.230072,0.231437,0.231635,0.234027,0.233746,0.236042,0.237874,0.237692,0.237647,0.237608,0.23757,0.237398,0.239075,0.239475,0.241573,0.241435,0.2414,0.241253,0.245604,0.245415,0.245241,0.247061,0.249642,0.252293,0.253826,0.253548,0.255771,0.255732,0.255554,0.257097,0.257805,0.257982,0.26083,0.2622,0.262028,0.262109,0.264953,0.26638,0.268053,0.268556,0.270461,0.267396,0.290604,0.290604,0.302114,0.302921,0.303762,0.30466,0.305635,0.30671,0.308051,0.309724,0.311495,0.313334,0.315211,0.317096,0.318959,0.320551,0.322033,0.323478,0.324895,0.326293,0.327684,0.329103,0.330574,0.332052,0.333537,0.335027,0.336522,0.338023,0.339601,0.34117,0.342719,0.344236,0.345709,0.347126,0.348331,0.349386,0.350411,0.35143,0.352469,0.353552,0.354773,0.356175,0.357661,0.359228,0.360877,0.362607,0.364431,0.36656,0.368732,0.370913,0.373067,0.375157,0.377149,0.378705,0.379751,0.380752,0.381778,0.382894,0.384168,0.385897,0.388629,0.391601,0.39475,0.398014,0.401331,0.40464,0.407803,0.410298,0.412702,0.415032,0.417309,0.41955,0.421774,0.424025,0.426318,0.428641,0.431006,0.433425,0.43591,0.438473,0.441273,0.444183,0.447166,0.450211,0.453308,0.456446,0.459612,0.462714,0.465834,0.468974,0.472134,0.475313,0.478512,0.481732,0.484977,0.488242,0.491526,0.494828,0.498148,0.501486,0.504836,0.508194,0.511569,0.514964,0.518381,0.52182,0.525282,0.528776,0.532303,0.535856,0.539433,0.543034,0.54666,0.550308,0.554043,0.557842,0.56164,0.565422,0.569174,0.572878,0.576522,0.579781,0.582868,0.585951,0.589074,0.59228,0.595612,0.599177,0.603669,0.608323,0.613083,0.617892,0.622691,0.627424,0.632033,0.635713,0.639235,0.642678,0.646087,0.649508,0.652984,0.656758,0.661055,0.665443,0.66989,0.674359,0.678819,0.683234,0.687267,0.690901,0.69452,0.698175,0.701915,0.705791,0.709854,0.715085,0.720672,0.726362,0.732065,0.737691,0.743153,0.748359,0.752328,0.755679,0.758831,0.76186,0.764842,0.767852,0.771296,0.775588,0.779951,0.784315,0.788607,0.792755,0.796688,0.799789,0.802379,0.80476,0.806978,0.809081,0.811118,0.813531,0.816236,0.81884,0.821278,0.823482,0.825384,0.826635,0.827013,0.827095,0.82695,0.826644,0.826247,0.826398,0.826784,0.827014,0.826994,0.826632,0.825834,0.823231,0.820269,0.817187,0.814173,0.811414,0.810308,0.810028,0.810045,0.810223,0.810421,0.810447,0.809372,0.808108,0.806699,0.805189,0.80362,0.802039,0.800489,0.799007,0.797635,0.796416,0.795415,0.794857,0.79453,0.794428,0.794547,0.794882,0.7955,0.796417,0.797496,0.798701,0.799997,0.801349,0.802723,0.804084,0.805392,0.806612,0.807706,0.80864,0.808934,0.808745,0.808515,0.808349,0.808351,0.808623,0.810127,0.812115,0.814391,0.81689,0.819544,0.822287,0.824613,0.826802,0.829044,0.831367,0.8338,0.836372,0.839311,0.842588,0.846008,0.849546,0.853175,0.856867,0.860549,0.863939,0.867372,0.870875,0.874475,0.878196,0.882065,0.8865,0.891238,0.896075,0.900961,0.905844,0.910675,0.915353,0.919418,0.923365,0.927219,0.931004,0.934744,0.938462,0.942157,0.945873,0.94965,0.953516,0.957501,0.961634,0.966224,0.971544,0.976954,0.982364,0.987684,0.992834,0.997704,1.001244,1.004074,1.006764,1.009424,1.012174,1.015134,1.019294,1.024644,1.030234,1.035944,1.041644,1.047194,1.052484,1.056524,1.060064,1.063264,1.066154,1.068744,1.071064,1.073044,1.074794,1.076374,1.077824,1.079184,1.080494,1.082214,1.083984,1.085674,1.087234,1.088614,1.089774,1.090464,1.090844,1.090934,1.090724,1.090204,1.089324,1.087854,1.086144,1.084234,1.082204,1.080104,1.078434,1.076884,1.075234,1.073414,1.071364,1.068724,1.064914,1.060994,1.057164,1.053594,1.050464,1.050014,1.050034,1.050264,1.050464,1.050384,1.049174,1.045904,1.042254,1.038394,1.034524,1.030924,1.028724,1.026814,1.025134,1.023604,1.022174,1.020764,1.019314,1.017774,1.016064,1.014144,1.011814,1.008424,1.004844,1.001214,0.997644,0.994274,0.992034,0.990154,0.988494,0.986994,0.985584,0.984204,0.982784,0.981284,0.979634,0.977794,0.975664,0.972224,0.968644,0.965104,0.961754,0.958781,0.957799,0.957748,0.957938,0.958146,0.958152,0.957635,0.955004,0.951916,0.948484,0.944823,0.941047,0.937493,0.934042,0.93071,0.927552,0.924624,0.9223,0.920475,0.918874,0.917437,0.916107,0.914825,0.913516,0.912146,0.910661,0.909006,0.907128,0.904299,0.900989,0.89766,0.894466,0.891565,0.889891,0.889726,0.889853,0.890066,0.890157,0.889919,0.887866,0.884916,0.881708,0.878398,0.875145,0.872638,0.87088,0.869345,0.867976,0.866719,0.865515,0.864299,0.863029,0.861652,0.860115,0.858365,0.855807,0.852649,0.849457,0.84638,0.843571,0.84171,0.841259,0.841173,0.84131,0.841524,0.841673,0.840974,0.839735,0.838327,0.836797,0.835188,0.833588,0.83217,0.830755,0.829341,0.827928,0.826516,0.825098,0.823679,0.822261,0.820845,0.819433,0.817966,0.81637,0.814833,0.813396,0.812102,0.810995,0.810848,0.811021,0.8112,0.811249,0.811032,0.810246,0.807614,0.804708,0.801706,0.798792,0.796144,0.795078,0.794657,0.794584,0.794769,0.795121,0.795476,0.795424,0.795372,0.795319,0.795266,0.795213,0.79526,0.795409,0.795497,0.795481,0.795322,0.794976,0.79406,0.792864,0.791513,0.790051,0.78852,0.786965,0.785431,0.783954,0.782575,0.781335,0.780276,0.779794,0.779576,0.779515,0.779571,0.779703,0.779836,0.779785,0.779735,0.779684,0.779633,0.779582,0.779531,0.77948,0.77943,0.779379,0.779328,0.779277,0.779224,0.779172,0.779119,0.779066,0.779014,0.778961,0.77891,0.778859,0.778808,0.778757,0.778706,0.778656,0.778605,0.778554,0.778503,0.778452,0.778401,0.77835,0.7783,0.778249,0.778198,0.778147,0.778096,0.778045,0.777994,0.777943,0.777892,0.777841,0.777791,0.77774,0.777689,0.777639,0.777588,0.777536,0.777484,0.777432,0.777379,0.777326,0.777273,0.777221,0.777169,0.777118,0.777067,0.777017,0.776966,0.776915,0.776865,0.776814,0.776763,0.776712,0.776661,0.77661,0.776559,0.776508,0.776457,0.776406,0.776356,0.776305,0.776254,0.776203,0.776152,0.776101,0.77605,0.775999,0.775948,0.775898,0.775847,0.775796,0.775745,0.775694,0.775643,0.775592,0.775541,0.77549,0.77544,0.775389,0.775338,0.775287,0.775236,0.775185,0.775134,0.775083,0.775032,0.774981,0.774931,0.77488,0.774829,0.774778,0.774727,0.774676,0.774625,0.774574,0.774523,0.774473,0.774422,0.774371,0.77432,0.774269,0.774218,0.774167,0.774116,0.774065,0.774014,0.773964,0.773913,0.773862,0.773811,0.77376,0.773817,0.773966,0.774055,0.774041,0.773884,0.773543,0.772488,0.771143,0.769722,0.768307,0.766981,0.766058,0.765748,0.765616,0.765621,0.765721,0.765877,0.765901,0.765852,0.765803,0.765754,0.765705,0.765655,0.765808,0.765929,0.76597,0.765893,0.765658,0.765056,0.763809,0.762445,0.761043,0.759684,0.758448,0.758066,0.758023,0.758066,0.758115,0.758089,0.75783,0.756624,0.755288,0.753901,0.752542,0.75129,0.750729,0.750663,0.750696,0.750749,0.750742,0.750595,0.749678,0.748529,0.747239,0.745847,0.744393,0.743001,0.741714,0.740429,0.739145,0.737864,0.73659,0.735543,0.734455,0.73328,0.731971,0.730481,0.728327,0.725624,0.722886,0.720244,0.717826,0.716171,0.715771,0.715687,0.715799,0.715982,0.716113,0.71555,0.714494,0.713292,0.711984,0.710607,0.709228,0.70801,0.706795,0.705581,0.704369,0.703159,0.701952,0.700748,0.699545,0.698343,0.697142,0.695904,0.694525,0.693192,0.691941,0.690812,0.689841,0.689671,0.689813,0.689967,0.690016,0.689844,0.689236,0.686993,0.684508,0.681937,0.679435,0.677155,0.676336,0.676121,0.676145,0.676293,0.67645,0.676412,0.675499,0.67443,0.673241,0.671966,0.670643,0.669305,0.66799,0.666734,0.665575,0.664547,0.663768,0.66347,0.663334,0.663323,0.6634,0.663531,0.663787,0.664106,0.664312,0.66433,0.664086,0.663505,0.661633,0.659281,0.656807,0.65436,0.65209,0.650765,0.650316,0.650178,0.650274,0.65053,0.650872,0.651046,0.651158,0.651207,0.651156,0.65097,0.650558,0.649655,0.648602,0.647434,0.646188,0.6449,0.643614,0.642359,0.641166,0.640069,0.639101,0.638432,0.638328,0.638333,0.63838,0.638401,0.638326,0.6377,0.636615,0.635451,0.634274,0.633153,0.632207,0.632077,0.632067,0.632111,0.632141,0.632088,0.631622,0.630569,0.629426,0.628258,0.627133,0.626117,0.625735,0.625564,0.625519,0.625568,0.625676,0.625744,0.625556,0.625403,0.625313,0.625315,0.625439,0.626161,0.627434,0.628686,0.629787,0.630604,0.631008,0.629978,0.627874,0.625519,0.623083,0.620742,0.619128,0.618634,0.618452,0.618512,0.618739,0.619063,0.619146,0.619106,0.619066,0.619025,0.618985,0.618945,0.618903,0.618861,0.618818,0.618776,0.618734,0.618692,0.618652,0.618612,0.618571,0.618531,0.618491,0.618449,0.618407,0.618365,0.618323,0.618281,0.618239,0.618198,0.618158,0.618117,0.618077,0.618037,0.617996,0.617954,0.617912,0.61787,0.617827,0.617785,0.61783,0.617948,0.618018,0.618007,0.617882,0.617611,0.616766,0.615692,0.614555,0.613422,0.612358,0.611589,0.611336,0.611225,0.611224,0.611301,0.611423,0.611448,0.611406,0.611364,0.611322,0.611279,0.611237,0.611196,0.611156,0.611116,0.611075,0.611035,0.610995,0.610955,0.610914,0.610874,0.610834,0.610793,0.610753,0.610713,0.610672,0.610632,0.610591,0.610551,0.610511,0.610471,0.610431,0.61039,0.61035,0.610309,0.610267,0.610225,0.610182,0.61014,0.610098,0.610056,0.610016,0.609975,0.609935,0.609895,0.609855,0.609815,0.609774,0.609734,0.609693,0.609653,0.609613,0.609572,0.609532,0.609492,0.609451,0.609411,0.609371,0.60933,0.60929,0.609249,0.609209,0.609169,0.609128,0.609088,0.609048,0.609007,0.608967,0.608927,0.608886,0.608846,0.608806,0.608766,0.608725,0.608648,0.608462,0.608312,0.608224,0.608227,0.60835,0.608876,0.609755,0.610713,0.611695,0.612645,0.613505,0.613929,0.614032,0.61402,0.613922,0.613765,0.613578,0.613527,0.613487,0.613447,0.613406,0.613366,0.613324,0.613282,0.61324,0.613198,0.613156,0.613114,0.613072,0.613032,0.612991,0.612951,0.612911,0.612871,0.612831,0.612791,0.61275,0.61271,0.612669,0.612628,0.612586,0.612544,0.612502,0.61246,0.612418,0.612376,0.612336,0.612295,0.612255,0.612215,0.612175,0.612134,0.612094,0.612054,0.612013,0.611973,0.611927,0.611739,0.61158,0.611479,0.611464,0.611563,0.611965,0.612824,0.613775,0.61476,0.615724,0.61661,0.617162,0.617292,0.617302,0.617219,0.617071,0.616887,0.616804,0.616762,0.616719,0.616677,0.616635,0.616593,0.616552,0.616512,0.616471,0.616431,0.616391,0.616351,0.616311,0.616271,0.61623,0.61619,0.616149,0.616012,0.615835,0.615705,0.615649,0.615697,0.615876,0.616655,0.617582,0.618567,0.619554,0.620485,0.621298,0.621485,0.621539,0.621488,0.621361,0.621186,0.620993,0.620811,0.620665,0.620585,0.620599,0.620734,0.621313,0.622208,0.623179,0.624171,0.625127,0.625991,0.626402,0.6265,0.626485,0.626383,0.626224,0.626034,0.62584,0.625673,0.625562,0.625537,0.625625,0.626296,0.628378,0.630291,0.631752,0.632475,0.632175,0.629457,0.623422,0.616874,0.610292,0.604154,0.60124,0.600076,0.599848,0.600361,0.601421,0.602754,0.603415,0.604209,0.605109,0.606088,0.607118,0.608053,0.608427,0.608913,0.609604,0.610596,0.611982,0.614408,0.61904,0.624085,0.629327,0.63455,0.639536,0.64407,0.647643,0.648515,0.648829,0.648707,0.64827,0.647641,0.647225,0.647181,0.647137,0.647093,0.647049,0.647006,0.646963,0.646921,0.646879,0.646837,0.646795,0.646753,0.646709,0.646665,0.646621,0.646577,0.646533,0.64649,0.646447,0.646405,0.646363,0.646321,0.646279,0.646136,0.645954,0.64582,0.645764,0.645817,0.646007,0.646826,0.647795,0.648824,0.649854,0.650826,0.651666,0.651705,0.651636,0.65152,0.651415,0.651379,0.651688,0.652598,0.653606,0.654652,0.655676,0.656618,0.657214,0.657354,0.657364,0.657276,0.65712,0.656924,0.656833,0.656789,0.656745,0.656701,0.656657,0.656612,0.65641,0.656238,0.656127,0.656107,0.656208,0.656565,0.657316,0.658205,0.659202,0.660278,0.661402,0.662547,0.663684,0.664781,0.665806,0.66673,0.667522,0.667991,0.668123,0.668127,0.668032,0.66787,0.66767,0.66759,0.667546,0.667502,0.667458,0.667414,0.66737,0.667327,0.667283,0.667239,0.667196,0.667151,0.66699,0.666663,0.666413,0.666299,0.666376,0.666701,0.668012,0.669909,0.671967,0.674071,0.676109,0.677967,0.679709,0.681191,0.68205,0.682111,0.681198;

bnd_Vol73 = 2.5813,2.5995,2.6178,2.63605,2.65431,2.67256,2.69081,2.70906,2.72731,2.74556,2.76381,2.78206,2.80032,2.8185,2.83682,2.85507,2.87332,2.89157,2.90982,2.92808,2.94633,2.96458,2.98283,3.00108,3.01933,3.03758,3.05584,3.07409,3.09234,3.11059,3.12884,3.14709,3.16534,3.18359,3.20185,3.2201,3.23835,3.2566,3.27485,3.2931,3.31135,3.32961,3.34786,3.36611,3.38436,3.40261,3.42086,3.43911,3.45736,3.47562,3.49387,3.51212,3.53037,3.54862,3.56687,3.58512,3.60338,3.62163,3.63988,3.65813,3.67638,3.69463,3.71288,3.73114,3.74939,3.76764,3.78589,3.80414,3.82239,3.84064,3.85889,3.87715,3.8954,3.91365,3.9319,3.95015,3.9684,3.98665,4.00491,4.02316,4.04141,4.05966,4.07791,4.09616,4.11441,4.13266,4.15092,4.16917,4.18742,4.20567,4.22392,4.24217,4.26042,4.27868,4.29693,4.31518,4.33343,4.35168,4.36993,4.38818,4.40643,4.42469,4.44294,4.46119,4.47944,4.49769,4.51594,4.53419,4.55245,4.5707,4.58895,4.6072,4.62545,4.6437,4.66195,4.68021,4.69846,4.71671,4.73496,4.75321,4.77146,4.78971,4.80796,4.82622,4.84447,4.86272,4.88097,4.89922,4.91747,4.93572,4.95398,4.97223,4.99048,5.00873,5.02698,5.04523,5.06348,5.08173,5.09999,5.11824,5.13649,5.15474,5.17299,5.19124,5.20949,5.22775,5.246,5.26425,5.2825,5.30075,5.319,5.33725,5.35551,5.37376,5.39201,5.41026,5.42851,5.44676,5.46501,5.48326,5.50152,5.51977,5.53802,5.55627,5.57452,5.59277,5.61102,5.62928,5.64753,5.66578,5.68403,5.70228,5.72053,5.73878,5.75703,5.77529,5.79354,5.81179,5.83004,5.84829,5.86654,5.88479,5.90305,5.9213,5.93955,5.9578,5.97605,5.9943,6.01255,6.03081,6.04906,6.06731,6.08556,6.10381,6.12206,6.14031,6.15856,6.17682,6.19507,6.21332,6.23157,6.24982,6.26807,6.28632,6.30458,6.32283,6.34108,6.35933,6.37758,6.39583,6.41408,6.43233,6.45059,6.46884,6.48709,6.50534,6.52359,6.54184,6.56009,6.57835,6.5966,6.61485,6.6331,6.65135,6.6696,6.68785,6.70611,6.72436,6.74261,6.76086,6.77911,6.79736,6.81561,6.83386,6.85212,6.87037,6.88862,6.90687,6.92512,6.94337,6.96162,6.97988,6.99813,7.01638,7.03463,7.05288,7.07113,7.08938,7.10763,7.12589,7.14414,7.16239,7.18064,7.19889,7.21714,7.23539,7.25365,7.2719,7.29015,7.3084,7.32665,7.3449,7.36315,7.38141,7.39966,7.41791,7.43616,7.45441,7.47266,7.49091,7.50916,7.52742,7.54567,7.56392,7.58217,7.60042,7.61867,7.63692,7.65518,7.67343,7.69168,7.70993,7.72818,7.74643,7.76468,7.78293,7.80119,7.81944,7.83769,7.85594,7.87419,7.89244,7.91069,7.92895,7.9472,7.96545,7.9837,8.00195,8.0202,8.03845,8.05671,8.07496,8.09321,8.11146,8.12971,8.14796,8.16621,8.18446,8.20272,8.22097,8.23922,8.25747,8.27572,8.29397,8.31222,8.33048,8.34873,8.36698,8.38523,8.40348,8.42173,8.43998,8.45823,8.47649,8.49474,8.51299,8.53124,8.54949,8.56774,8.58599,8.60425,8.6225,8.64075,8.659,8.67725,8.6955,8.71375,8.732,8.75026,8.76851,8.78676,8.80501,8.82326,8.84151,8.85976,8.87802,8.89627,8.91452,8.93277,8.95102,8.96927,8.98752,9.00578,9.02403,9.04228,9.06053,9.07878,9.09703,9.11528,9.13353,9.15179,9.17004,9.18829,9.20654,9.22479,9.24304,9.26129,9.27955,9.2978,9.31605,9.3343,9.35255,9.3708,9.38905,9.4073,9.42556,9.44381,9.46206,9.48031,9.49856,9.51681,9.53506,9.55332,9.57157,9.58982,9.60807,9.62632,9.64457,9.66282,9.68108,9.69933,9.71758,9.73583,9.75408,9.77233,9.79058,9.80883,9.82709,9.84534,9.86359,9.88184,9.90009,9.91834,9.93659,9.95485,9.9731,9.99135,10.0096,10.0279,10.0461,10.0644,10.0826,10.1009,10.1191,10.1374,10.1556,10.1739,10.1921,10.2104,10.2286,10.2469,10.2651,10.2834,10.3016,10.3199,10.3381,10.3564,10.3746,10.3929,10.4111,10.4294,10.4476,10.4659,10.4841,10.5024,10.5206,10.5389,10.5571,10.5754,10.5936,10.6119,10.6301,10.6484,10.6666,10.6849,10.7032,10.7214,10.7397,10.7579,10.7762,10.7944,10.8127,10.8309,10.8492,10.8674,10.8857,10.9039,10.9222,10.9404,10.9587,10.9769,10.9952,11.0134,11.0317,11.0499,11.0682,11.0864,11.1047,11.1229,11.1412,11.1594,11.1777,11.1959,11.2142,11.2324,11.2507,11.2689,11.2872,11.3054,11.3237,11.3419,11.3602,11.3785,11.3967,11.415,11.4332,11.4515,11.4697,11.488,11.5062,11.5245,11.5427,11.561,11.5792,11.5975,11.6157,11.634,11.6522    ,11.6705,11.6887,11.707,11.7252,11.7435,11.7617,11.78,11.7982,11.8165,11.8347,11.853,11.8712,11.8895,11.9077,11.926,11.9442,11.9625,11.9807,11.999,12.0172,12.0355,12.0538,12.072,12.0903,12.1085,12.1268,12.145,12.1633,12.1815,12.1998,12.218,12.2363,12.2545,12.2728,12.291,12.3093,12.3275,12.3458,12.364,12.3823,12.4005,12.4188,12.437,12.4553,12.4735,12.4918,12.51,12.5283,12.5465,12.5648,12.583,12.6013,12.6195,12.6378,12.656,12.6743,12.6925,12.7108,12.7291,12.7473,12.7656,12.7838,12.8021,12.8203,12.8386,12.8568,12.8751,12.8933,12.9116,12.9298,12.9481,12.9663,12.9846,13.0028,13.0211,13.0393,13.0576,13.0758,13.0941,13.1123,13.1306,13.1488,13.1671,13.1853,13.2036,13.2218,13.2401,13.2583,13.2766,13.2948,13.3131,13.3313,13.3496,13.3678,13.3861,13.4044,13.4226,13.4409,13.4591,13.4774,13.4956,13.5139,13.5321,13.5504,13.5686,13.5869,13.6051,13.6234,13.6416,13.6599,13.6781,13.6964,13.7146,13.7329,13.7511,13.7694,13.7876,13.8059,13.8241,13.8424,13.8606,13.8789,13.8971,13.9154,13.9336,13.9519,13.9701,13.9884,14.0066,14.0249,14.0431,14.0614,14.0797,14.0979,14.1162,14.1344,14.1527,14.1709,14.1892,14.2074,14.2257,14.2439,14.2622,14.2804,14.2987,14.3169,14.3352,14.3534,14.3717,14.3899,14.4082,14.4264,14.4447,14.4629,14.4812,14.4994,14.5177,14.5359,14.5542,14.5724,14.5907,14.6089,14.6272,14.6454,14.6637,14.6819,14.7002,14.7184,14.7367,14.755,14.7732,14.7915,14.8097,14.828,14.8462,14.8645,14.8827,14.901,14.9192,14.9375,14.9557,14.974,14.9922,15.0105,15.047,15.0652,15.0835,15.12,15.1382,15.1565,15.1747,15.193,15.2112,15.2295,15.2477,15.266,15.2842,15.3025,15.3207,15.339,15.3572,15.3755,15.3937,15.412,15.4303,15.4485,15.4668,15.485,15.5033,15.5215,15.5398,15.558,15.5763,15.5945,15.6128,15.631,15.6493,15.6675,15.6858,15.704,15.7223,15.7405,15.7588,15.777,15.7953,15.8135,15.8318,15.85,15.8683,15.8865,15.9048,15.923,15.9413,15.9595,15.9778,15.996,16.0143,16.1421,16.1603,16.1786,16.1968,16.2151,16.2333,16.2516,16.2698,16.2881,16.3063,16.3246,16.3428,16.3611,16.3793,16.3976,16.4158,16.4341,16.4523,16.4706,16.4888,16.5071,16.5253,16.5436,16.5618,16.5801,16.5983,16.6166,16.6348,16.6531,16.6713,16.6896,16.7078,16.7261,16.7443,16.7626,16.7809,16.7991,16.8174,16.8356,16.8539,16.8721,16.8904,16.9086,16.9269,16.9451,16.9634,16.9816,16.9999,17.0181,17.0364,17.0546,17.0729,17.0911,17.1094,17.1276,17.1459,17.1641,17.1824,17.2006,17.2189,17.2371,17.2554,17.2736,17.2919,17.3101,17.3284,17.3466,17.3649,17.3831,17.4014,17.4196,17.4379,17.4562,17.4744,17.4927,17.5109,17.5292,17.5474,17.5657,17.5839,17.6022,17.6204,17.6387,17.6569,17.6752,17.6934,17.7117,17.7299,17.7482,17.7664,17.7847,17.8029,17.8212,17.8394,17.8577,17.8759,17.8942,17.9124,17.9307,17.9489,17.9672,17.9854,18.0037,18.0219,18.0402,18.0584,18.0767,18.0949,18.1132,18.1315,18.1497,18.168,18.1862,18.2045,18.2227,18.241,18.2592,18.2775,18.2957,18.314,18.3322,18.3505,18.3687,18.387,18.4052,18.4235,18.4417,18.46,18.4782,18.4965,18.5147,18.533,18.5512,18.5695,18.5877,18.606,18.6242,18.6425,18.6607,18.679,18.6972,18.7155,18.7337,18.752,18.7702,18.7885,18.8068,18.825,18.8433,18.8615,18.8798,18.898,18.9163,18.9345,18.9528,18.971,18.9893,19.0075,19.0258,19.044,19.0623,19.0805,19.0988,19.117,19.1353,19.1535,19.1718,19.19,19.2083,19.2265,19.2448,19.263,19.2813,19.2995,19.3178,19.336,19.3543,19.3725,19.3908,19.409,19.4273,19.4455,19.4638,19.4821,19.5003,19.5186,19.5368,19.5551,19.5733,19.5916,19.6098,19.6281,19.6463,19.6646,19.6828,19.7011,19.7193,19.7376,19.7558,19.7741,19.7923,19.8106,19.8288,19.8471,19.8653,19.8836,19.9018,19.9201,19.9383,19.9566,19.9748,19.9931,20.0113,20.0296,20.0478,20.0661,20.0843,20.1026,20.1208,20.1391,20.1574,20.1756,20.1939,20.2121,20.2304,20.2486,20.2669,20.2851,20.3034,20.3216,20.3399,20.3581,20.3764,20.3946,20.4129,20.4311,20.4494,20.4676,20.4859,20.5041,20.5224,20.5406,20.5589,20.5771,20.5954,20.6136,20.6319,20.6501,20.6684,20.6866,20.7049,20.7231,20.7414,20.7596,20.7779,20.7961,20.8144,20.8326,20.8509,20.8692,20.8874,20.9057,20.9239,20.9422,20.9604,20.9787,20.9969,21.0152,21.0334,21.0517,21.0699,21.0882,21.1064,21.1247,21.1429,21.1612,21.1794,21.1977,21.2159,21.2342,21.2524,21.2707,21.2889,21.3072,21.3254,21.3437,21.3619,21.3802,21.3984,21.4167,21.4349,21.4532,21.4714,21.4897,21.5079,21.5262,21.5445,21.5627,21.581,21.5992,21.6175,21.6357,21.654,21.6722,21.6905,21.7087,21.727,21.7452,21.7635,21.7817,21.8,21.8182,21.8365,21.8547,21.873,21.8912,21.9095,21.9277,21.946,21.9642,21.9825,22.0007,22.019,22.0372,22.0555,22.0737,22.092,22.1102,22.1285,22.1467,22.165,22.1832,22.2015,22.2198,22.238,22.2563,22.2745,22.2928,22.311,22.3293,22.3475,22.3658,22.384,22.4023,22.4205,22.4388,22.457,22.4753,22.4935,22.5118,22.53,22.5483,22.5665,22.5848,22.603,22.6213,22.6395,22.6578,22.676,22.6943,22.7125,22.7308,22.749,22.7673,22.7855,22.8038,22.822,22.8403,22.8585,22.8768,22.8951,22.9133,22.9316,22.9498,22.9681,22.9863,23.0046,23.0228,23.0411,23.0593,23.0776,23.0958,23.1141,23.1323,23.1506,23.1688,23.1871,23.2053,23.2236,23.2418,23.2601,23.2783,23.2966,23.3148,23.3331,23.3513,23.3696,23.3878,23.4061,23.4243,23.4426,23.4608,23.4791,23.4973,23.5156,23.5338,23.5521,23.5704,23.5886,23.6069,23.6251,23.6434,23.6616,23.6799,23.6981,23.7164,23.7346,23.7529,23.7711,23.7894,23.8076,23.8259,23.8441,23.8624,23.8806,23.8989,23.9171,23.9354,23.9536,23.9719,23.9901,24.0084,24.0266,24.0449,24.0631,24.0814,24.0996,24.1179,24.1361,24.1544,24.1726,24.1909,24.2091,24.2274,24.2457,24.2639,24.2822,24.3004,24.3187,24.3369,24.3552,24.3734,24.3917,24.4099,24.4282,24.4464,24.4647,24.4829,24.5012,24.5194,24.5377,24.5559,24.5742,24.5924,24.6107,24.6289,24.6472,24.6654,24.6837,24.7019,24.7202,24.7384,24.7567,24.7749,24.7932,24.8114,24.8297,24.8479,24.8662,24.8844,24.9027,24.921,24.9392,24.9575,24.9757,24.994,25.0122,25.0305,25.0487,25.067,25.0852,25.1035,25.1217,25.14,25.1582,25.1765,25.1947,25.213,25.2312,25.2495,25.2677,25.286,25.3042,25.3225,25.3407,25.359,25.3772,25.3955,25.4137,25.432,25.4502,25.4685,25.4867,25.505,25.5232,25.5415,25.5597,25.578,25.5963,25.6145,25.6328,25.651,25.6693,25.6875,25.7058,25.724,25.7423,25.7605,25.7788,25.797,25.8153,25.8335,25.8518,25.87,25.8883,25.9065,25.9248,25.943,25.9613,25.9795,25.9978,26.016,26.0343,26.0525,26.0708,26.089,26.1073,26.1255,26.1438,26.162,26.1803,26.1985,26.2168,26.235,26.2533,26.2716,26.2898,26.3081,26.3263,26.3446,26.3628,26.3811,26.3993,26.4176,26.4358,26.4541,26.4723,26.4906,26.5088,26.5271,26.5453,26.5636,26.5818,26.6001,26.6183,26.6366,26.6548,26.6731,26.6913,26.7096,26.7278,26.7461,26.7643,26.7826,26.8008,26.8191,26.8373,26.8556,26.8738,26.8921,26.9103,26.9286,26.9469,26.9651,26.9834,27.0016,27.0199,27.0381,27.0564,27.0746,27.0929,27.1111,27.1294,27.1476,27.1659,27.1841,27.2024,27.2206,27.2389,27.2571,27.2754,27.2936,27.3119,27.3301,27.3484,27.3666,27.3849,27.4031,27.4214,27.4396,27.4579,27.4761,27.4944,27.5126,27.5309,27.5491,27.5674,27.5856,27.6039,27.6222,27.6404,27.6587,27.6769,27.6952,27.7134,27.7317,27.7499,27.7682,27.7864,27.8047,27.8229,27.8412,27.8594,27.8777,27.8959,27.9142,27.9324,27.9507,27.9689,27.9872,28.0054,28.0237,28.0419,28.0602,28.0784,28.0967,28.1149,28.1332,28.1514,28.1697,28.1879,28.2062,28.2244,28.2427,28.2609,28.2792,28.2975,28.3157,28.334,28.3522,28.3705,28.3887,28.407,28.4252,28.4435,28.4617,28.48,28.4982,28.5165,28.5347,28.553,28.5712,28.5895,28.6077,28.626,28.6442,28.6625,28.6807,28.699,28.7172,28.7355,28.7537,28.772,28.7902,28.8085,28.8267,28.845,28.8632,28.8815,28.8997,28.918,28.9362,28.9545,28.9728,28.991,29.0093,29.0275,29.0458,29.064,29.0823,29.1005,29.1188,29.137,29.1553,29.1735,29.1918,29.21,29.2283,29.2465,29.2648,29.283,29.3013,29.3195,29.3378,29.356,29.3743,29.3925,29.4108,29.429,29.4473,29.4655,29.4838,29.502,29.5203,29.5385,29.5568,29.575,29.5933,29.6115,29.6298,29.6481,29.6663,29.6846,29.7028,29.7211,29.7393,29.7576,29.7758,29.7941,29.8123,29.8306,29.8488,29.8671,29.8853,29.9036,29.9218,29.9401,29.9583,29.9766,29.9948,30.0131,30.0313,30.0496,30.0678,30.0861,30.1043,30.1226,30.1408,30.1591,30.1773,30.1956,30.2138,30.2321,30.2503,30.2686,30.2868,30.3051,30.3234,30.3416,30.3599,30.3781,30.3964,30.4146,30.4329,30.4511,30.4694,30.4876,30.5059,30.5241,30.5424,30.5606,30.5789,30.5971,30.6154,30.6336,30.6519,30.6701,30.6884,30.7066,30.7249,30.7431,30.7614,30.7796,30.7979,30.8161,30.8344,30.8526,30.8709,30.8891,30.9074,30.9256,30.9439,30.9621,30.9804,30.9987,31.0169,31.0352,31.0534,31.0717,31.0899,31.1082,31.1264,31.1447,31.1629,31.1812,31.1994,31.2177,31.2359,31.2542,31.2724,31.2907,31.3089,31.3272,31.3454,31.3637,31.3819,31.4002,31.4184,31.4367,31.4549,31.4732,31.4914,31.5097,31.5279,31.5462,31.5644,31.5827,31.6009,31.6192,31.6374,31.6557,31.674,31.6922,31.7105,31.7287,31.747,31.7652,31.7835,31.8017,31.82,31.8382,31.8565,31.8747,31.893,31.9112,31.9295,31.9477,31.966,31.9842,32.0025,32.0207,32.039,32.0572,32.0755,32.0937,32.112,32.1302,32.1485,32.1667,32.185,32.2032,32.2215,32.2397,32.258,32.2762,32.2945,32.3127,32.331,32.3493,32.3675,32.3858,32.404,32.4223,32.4405,32.4588,32.477,32.4953,32.5135,32.5318,32.55,32.5683,32.5865,32.6048,32.623,32.6413,32.6595,32.6778,32.696,32.7143,32.7325,32.7508,32.769,32.7873,32.8055,32.8238,32.842,32.8603,32.8785,32.8968,32.915,32.9333,32.9515,32.9698,32.988,33.0063,33.0246,33.0428,33.0611,33.0793,33.0976,33.1158,33.1341,33.1523,33.1706,33.1888,33.2071,33.2253,33.2436,33.2618,33.2801,33.2983,33.3166,33.3348,33.3531,33.3713,33.3896,33.4078,33.4261,33.4443,33.4626,33.4808,33.4991,33.5173,33.5356,33.5538,33.5721,33.5903,33.6086,33.6268,33.6451,33.6633,33.6816,33.6999,33.7181,33.7364,33.7546,33.7729,33.7911,33.8094,33.8276,33.8459,33.8641,33.8824,33.9006,33.9189,33.9371,33.9554,33.9736,33.9919,34.0101,34.0284,34.0466,34.0649,34.0831,34.1014,34.1196,34.1379,34.1561,34.1744,34.1926,34.2109,34.2291,34.2474,34.2656,34.2839,34.3021,34.3204,34.3386,34.3569,34.3752,34.3934,34.4117,34.4299,34.4482,34.4664,34.4847,34.5029,34.5212,34.5394,34.5577,34.5759,34.5942,34.6124,34.6307,34.6489,34.6672,34.6854,34.7037,34.7219,34.7402,34.7584,34.7767,34.7949,34.8132,34.8314,34.8497,34.8679,34.8862,34.9044,34.9227,34.9409,34.9592,34.9774,34.9957,35.0139,35.0322,35.0505,35.0687,35.087,35.1052,35.1235,35.1417,35.16,35.1782,35.1965,35.2147,35.233,35.2512,35.2695,35.2877,35.306,35.3242,35.3425,35.3607,35.379,35.3972,35.4155,35.4337,35.452,35.4702,35.4885,35.5067,35.525,35.5432,35.5615,35.5797,35.598,35.6162,35.6345,35.6527,35.671,35.6892,35.7075,35.7258,35.744,35.7623,35.7805,35.7988,35.817,35.8353,35.8535,35.8718,35.89,35.9083,35.9265,35.9448,35.963,35.9813,35.9995,36.0178,36.036,36.0543,36.0725,36.0908,36.109,36.1273,36.1455,36.1638,36.182,36.2003,36.2185,36.2368,36.255,36.2733,36.2915,36.3098,36.328,36.3463,36.3645,36.3828,36.4011,36.4193,36.4376,36.4558,36.4741,36.4923,36.5106,36.5288,36.5471,36.5653,36.5836,36.6018,36.6201,36.6383,36.6566,36.6748,36.6931,36.7113,36.7296,36.7478,36.7661,36.7843,36.8026,36.8208,36.8391,36.8573,36.8756,36.8938,36.9121,36.9303,36.9486,36.9668,36.9851,37.0033,37.0216,37.0398,37.0581,37.0764,37.0946,37.1129,37.1311,37.1494,37.1676,37.1859,37.2041,37.2224,37.2406,37.2589,37.2771,37.2954,37.3136,37.3319,37.3501,37.3684,37.3866,37.4049,37.4231,37.4414,37.4596,37.4779,37.4961,37.5144,37.5326,37.5509,37.5691,37.5874,37.6056,37.6239,37.6421,37.6604,37.6786,37.6969,37.7151,37.7334,37.7517,37.7699,37.7882,37.8064,37.8247,37.8429,37.8612,37.8794,37.8977,37.9159,37.9342,37.9524,37.9707,37.9889,38.0072,38.0254,38.0437,38.0619,38.0802,38.0984,38.1167,38.1349,38.1532,38.1714,38.1897,38.2079,38.2262,38.2444,38.2627,38.2809,38.2992,38.3174,38.3357,38.3539,38.3722,38.3904,38.4087,38.427,38.4452,38.4635,38.4817,38.5,38.5182,38.5365,38.5547,38.573,38.5912,38.6095,38.6277,38.646,38.6642,38.6825,38.7007,38.719,38.7372,38.7555,38.7737,38.792,38.8102,38.8285,38.8467,38.865,38.8832,38.9015,38.9197,38.938,38.9562,38.9745,38.9927,39.011,39.0292,39.0475,39.0657,39.084;
idx_rfr_Vol73_rl = 1.4529,1.45264,1.45237,1.45207,1.45626,1.45554,1.45918,1.45947,1.45896,1.4623,1.46321,1.46707,1.46656,1.4663,1.46584,1.4685,1.46974,1.46815,1.46764,1.46487,1.46447,1.46428,1.46401,1.46375,1.46324,1.4669,1.46781,1.47113,1.47373,1.4789,1.48111,1.48696,1.49003,1.4951,1.50041,1.50264,1.5022,1.50193,1.50167,1.50144,1.49531,1.49293,1.48329,1.47715,1.4754,1.46632,1.46075,1.4576,1.45715,1.45972,1.46106,1.4606,1.4628,1.46453,1.46416,1.46395,1.46374,1.46338,1.46505,1.4671,1.47102,1.47076,1.47057,1.4703,1.47004,1.46977,1.46946,1.47366,1.47294,1.47675,1.47317,1.47685,1.47634,1.47607,1.47581,1.47554,1.47522,1.47676,1.47913,1.47878,1.48287,1.48237,1.48211,1.48179,1.48405,1.4856,1.48537,1.48486,1.48821,1.48878,1.48851,1.48825,1.48798,1.48772,1.48745,1.48719,1.48692,1.48666,1.4864,1.48624,1.48596,1.4857,1.48525,1.48781,1.48916,1.48977,1.49303,1.49225,1.50076,1.50031,1.49991,1.50401,1.50373,1.5033,1.50718,1.50715,1.5067,1.51032,1.51056,1.51035,1.51014,1.51038,1.514,1.51355,1.51352,1.5172,1.51968,1.52078,1.52481,1.52676,1.52837,1.53293,1.53617,1.54167,1.54406,1.55238,1.5559,1.55994,1.56808,1.5741,1.58222,1.59016,1.5963,1.60056,1.60009,1.60011,1.58901,1.56809,1.55453,1.54222,1.52777,1.50799,1.49571,1.48926,1.48046,1.47441,1.46841,1.46313,1.45835,1.45405,1.45308,1.44962,1.4453,1.44503,1.44198,1.44023,1.43545,1.43547,1.43521,1.43514,1.43198,1.43029,1.43004,1.42977,1.42951,1.42925,1.42898,1.42862,1.43299,1.43012,1.42783,1.43214,1.4317,1.43144,1.43061,1.42641,1.42627,1.4305,1.43037,1.42655,1.42548,1.42521,1.42495,1.42468,1.42467,1.42094,1.41978,1.41952,1.41925,1.41899,1.41872,1.41846,1.41819,1.41796,1.41777,1.4175,1.41724,1.41697,1.4167,1.41644,1.41618,1.41591,1.41564,1.41544,1.41522,1.41495,1.41469,1.41442,1.41416,1.41389,1.41363,1.41336,1.41315,1.41294,1.41315,1.4168,1.41636,1.41605,1.41733,1.41996,1.4195,1.42042,1.42316,1.42656,1.42678,1.42636,1.42951,1.43447,1.4339,1.43683,1.4378,1.43878,1.44145,1.44501,1.44592,1.44935,1.44866,1.45288,1.45252,1.45225,1.45199,1.45172,1.45146,1.4512,1.45093,1.45073,1.45052,1.44734,1.44731,1.4455,1.4393,1.43647,1.43589,1.42746,1.42416,1.41807,1.41197,1.40599,1.39995,1.39419,1.38411,1.37971,1.37142,1.36421,1.35125,1.34861,1.33862,1.32821,1.32032,1.31529,1.30477,1.29506,1.28935,1.27672,1.26835,1.26168,1.24882,1.24176,1.23324,1.22917,1.21764,1.20862,1.20232,1.19461,1.18663,1.18376,1.17407,1.16845,1.16682,1.16056,1.15451,1.14852,1.14243,1.13645,1.13036,1.12438,1.1181,1.11617,1.106,1.09999,1.09844,1.08912,1.09005,1.08069,1.07905,1.07261,1.07188,1.06969,1.06331,1.06184,1.05821,1.05397,1.05355,1.05358,1.04902,1.04839,1.05068,1.05231,1.05174,1.05511,1.06559,1.07536,1.09329,1.11348,1.14597,1.17689,1.22532,1.30264,1.38057,1.42693,1.45127,1.49094,1.55463,1.54141,1.59183,1.70822,1.76198,1.77635,1.81618,1.83904,1.84817,1.85324,1.8596,1.87458,1.89342,1.91532,1.93429,1.95349,1.99517,2.07046,2.13625,2.16891,2.2063,2.23525,2.30465,2.37685,2.43263,2.48099,2.527,2.57085,2.61661,2.66245,2.70069,2.74143,2.77705,2.80653,2.84703,2.88426,2.90868,2.92736,2.95346,2.97869,2.99297,3.00569,3.01564,3.02178,3.02604,3.02594,3.02173,3.01456,3.00178,2.99397,2.97041,2.95516,2.93153,2.91683,2.88861,2.86172,2.82834,2.79689,2.76196,2.73776,2.70735,2.68009,2.65252,2.61922,2.5926,2.56153,2.5302,2.5061,2.47724,2.45778,2.42248,2.39074,2.36638,2.33483,2.29458,2.25206,2.21814,2.17314,2.13909,2.10185,2.07171,2.04827,2.03271,2.00855,1.98192,1.94813,1.92771,1.88735,1.8504,1.81442,1.78302,1.77478,1.75021,1.73177,1.71934,1.71271,1.70681,1.70068,1.69914,1.69562,1.69561,1.69617,1.70347,1.71385,1.71987,1.73057,1.7436,1.75324,1.76318,1.77306,1.78301,1.79316,1.80032,1.80547,1.81367,1.81271,1.81637,1.821,1.82061,1.82016,1.82444,1.82839,1.82787,1.8277,1.82744,1.82788,1.81827,1.81833,1.81807,1.81784,1.81303,1.81327,1.80865,1.80842,1.80816,1.8079,1.80763,1.80736,1.8071,1.80687,1.80667,1.8064,1.80614,1.80588,1.80561,1.80535,1.80509,1.80483,1.80361,1.79997,1.79991,1.79965,1.79969,1.79538,1.79475,1.79448,1.79422,1.79409,1.79127,1.78917,1.78906,1.78879,1.78871,1.78381,1.78378,1.78352,1.78328,1.7831,1.78282,1.78256,1.7826,1.77834,1.77758,1.7774,1.77713,1.7762,1.7721,1.77213,1.77196,1.76947,1.76715,1.76711,1.76441,1.76222,1.76206,1.7618,1.76171,1.7568,1.75709,1.75276,1.75216,1.7519,1.75162,1.75054,1.74671,1.74672,1.74571,1.7417,1.74173,1.74056,1.73687,1.73682,1.73656,1.7363,1.73602,1.73576,1.73549,1.73532,1.73506,1.73454,1.73813,1.73417,1.73401,1.73375,1.73376,1.73769,1.73716,1.73689,1.73662,1.73643,1.73621,1.73593,1.73567,1.73541,1.73515,1.73487,1.73461,1.73435,1.73408,1.73403,1.72916,1.72949,1.72482,1.72475,1.72163,1.71984,1.71507,1.71548,1.71069,1.70889,1.70896,1.70567,1.70715,1.70685,1.70498,1.70473,1.70447,1.70421,1.70394,1.70367,1.70351,1.70325,1.70298,1.70272,1.70246,1.7025,1.69812,1.6967,1.69281,1.69281,1.69146,1.68823,1.68369,1.68366,1.68065,1.6745,1.67433,1.67436,1.66946,1.66491,1.66523,1.66052,1.65852,1.65568,1.65513,1.64891,1.64661,1.64581,1.6395,1.63754,1.63754,1.63473,1.62868,1.62846,1.62513,1.62351,1.61883,1.61887,1.6186,1.61734,1.61077,1.60952,1.60776,1.6049,1.60027,1.60033,1.59682,1.5911,1.59101,1.59074,1.59009,1.58361,1.58152,1.58137,1.58139,1.57733,1.57657,1.57395,1.57166,1.57059,1.56712,1.56277,1.56235,1.56209,1.56182,1.5607,1.55697,1.55702,1.55218,1.55228,1.55215,1.54727,1.5475,1.54304,1.54263,1.54237,1.5422,1.53757,1.53457,1.533,1.53292,1.52957,1.52781,1.52339,1.52389,1.5145,1.51451,1.51471,1.50379,1.48724,1.48884,1.50575,1.51041,1.51373,1.50917,1.49868,1.49776,1.49687,1.49603,1.49526,1.49459,1.49431,1.49441,1.49454,1.49461,1.49456,1.49431,1.49312,1.49149,1.48976,1.48804,1.48644,1.48542,1.48519,1.48515,1.48522,1.48533,1.4854,1.48501,1.48434,1.48358,1.48275,1.48187,1.48097,1.48007,1.47918,1.47835,1.47759,1.47693,1.47654,1.47638,1.47631,1.47633,1.47639,1.47648,1.47672,1.47693,1.47706,1.47703,1.47681,1.47626,1.47475,1.47307,1.46718,1.46738,1.4676,1.46758,1.46756,1.46755,1.46753,1.46751,1.46749,1.46746,1.46743,1.46739,1.46735,1.46732,1.46721,1.46708,1.46698,1.46693,1.46695,1.46707,1.46759,1.46826,1.46898,1.46971,1.4704,1.47102,1.47113,1.47109,1.471,1.47092,1.47087,1.47093,1.47133,1.47184,1.47246,1.47321,1.47406,1.47506,1.47634,1.47769,1.47908,1.48046,1.48181,1.48309,1.48345,1.4838,1.48426,1.48491,1.48587,1.48726,1.49074,1.49472,1.49909,1.50373,1.50854,1.51341,1.51822,1.52196,1.52473,1.52747,1.53028,1.53326,1.5365,1.54011,1.54582,1.55274,1.56016,1.56796,1.57605,1.58432,1.59265,1.60095,1.6091,1.617,1.62454,1.63161,1.63811,1.64394,1.64897,1.65312,1.65626,1.65953,1.67091,1.68322,1.69635,1.71016,1.72455,1.73939,1.75456,1.76995,1.78543,1.80089,1.8162,1.83125,1.84592,1.86008,1.87363,1.88643,1.89837,1.90933,1.9192,1.92296,1.92533,1.92826,1.93172,1.93567,1.94008,1.94491,1.95013,1.95571,1.9616,1.96777,1.97419,1.98083,1.98764,1.9946,2.0017,2.00916,2.01663,2.02405,2.03137,2.03851,2.04542,2.05204,2.05831,2.0637,2.06581,2.06798,2.07045,2.07352,2.07743,2.08246,2.08948,2.10664,2.1256,2.14584,2.16686,2.18817,2.20925,2.22961,2.24874,2.26614,2.27899,2.28481,2.28902,2.2918,2.29336,2.29388,2.29355,2.29294,2.29193,2.29043,2.28853,2.28631,2.28404,2.28185,2.27949,2.27694,2.27421,2.27118,2.26773,2.26418,2.26062,2.25713,2.25405,2.25153,2.2491,2.24669,2.24421,2.24135,2.23779,2.2342,2.23066,2.2273,2.22456,2.22259,2.2209,2.2194,2.21805,2.21669,2.21486,2.21308,2.21142,2.20992,2.20863,2.20812,2.20797,2.20798,2.20807,2.20817,2.20816,2.20732,2.20642,2.20553,2.20471,2.20405,2.20387,2.20419,2.20474,2.20548,2.20639,2.20744,2.20857,2.20976,2.21103,2.21237,2.21374,2.21515,2.21646,2.2176,2.2188,2.22006,2.22142,2.22291,2.22469,2.2271,2.22963,2.23223,2.23483,2.23738,2.23982,2.24165,2.24301,2.24429,2.24554,2.24682,2.24818,2.24991,2.25208,2.25442,2.2569,2.25952,2.26224,2.26507,2.26794,2.27087,2.27386,2.2769,2.27997,2.28307,2.28619,2.28894,2.29173,2.2946,2.29759,2.30075,2.30412,2.30789,2.31264,2.31765,2.32286,2.32821,2.33366,2.33914,2.34462,2.34985,2.35444,2.35895,2.36341,2.36784,2.37225,2.37666,2.3811,2.38577,2.39055,2.39537,2.40022,2.4051,2.41,2.41492,2.41985,2.4248,2.42976,2.43469,2.43961,2.4445,2.44935,2.45415,2.45884,2.46337,2.46786,2.47231,2.47672,2.48111,2.48548,2.48985,2.49441,2.49898,2.50352,2.50802,2.51245,2.51681,2.52106,2.52501,2.52851,2.53197,2.53542,2.53891,2.54249,2.54621,2.55037,2.55523,2.56028,2.56549,2.5708,2.5762,2.58164,2.58709,2.59219,2.5968,2.60143,2.60612,2.61092,2.61586,2.62099,2.62635,2.63299,2.64027,2.64778,2.65545,2.66321,2.671,2.67875,2.68638,2.69383,2.70082,2.70707,2.71302,2.71867,2.72401,2.72902,2.73368,2.73798,2.74158,2.74432,2.74684,2.74924,2.7516,2.75401,2.75655,2.7599,2.76367,2.76771,2.77202,2.7766,2.78146,2.78659,2.79216,2.79844,2.80495,2.81162,2.81841,2.82527,2.83213,2.83894,2.84565,2.85178,2.85736,2.86281,2.86812,2.87333,2.87843,2.88346,2.88842,2.89358,2.89886,2.90405,2.90911,2.91403,2.91877,2.92331,2.92761,2.93109,2.9343,2.93736,2.94031,2.9432,2.94607,2.949,2.95241,2.95589,2.95943,2.963,2.96661,2.97023,2.97386,2.97749,2.9811,2.98469,2.98825,2.99177,2.99523,2.99862,3.00178,3.00486,3.0079,3.0109,3.01387,3.01683,3.0198,3.02295,3.02609,3.0292,3.03228,3.03531,3.03827,3.04116,3.04396,3.04666,3.04924,3.05168,3.05398,3.05611,3.05802,3.05973,3.06124,3.06255,3.06366,3.06455,3.06508,3.06528,3.06533,3.06524,3.06508,3.06486,3.06478,3.06474,3.06471,3.06467,3.06464,3.0646,3.06457,3.06453,3.0645,3.06446,3.06443,3.06446,3.06469,3.06485,3.06489,3.06477,3.06443,3.06354,3.06218,3.06061,3.0589,3.0571,3.05535,3.05387,3.05236,3.05077,3.04907,3.04724,3.04485,3.04233,3.03977,3.03724,3.0348,3.033,3.03142,3.02989,3.02835,3.02673,3.02473,3.02235,3.01985,3.01727,3.01464,3.0122,3.01003,3.00774,3.00526,3.00248,2.99905,2.9947,2.99011,2.98544,2.98081,2.97679,2.97319,2.96974,2.96638,2.96308,2.95942,2.95571,2.95212,2.94875,2.94565,2.94376,2.94221,2.94077,2.9393,2.93764,2.9351,2.93187,2.9284,2.92476,2.92103,2.91739,2.91382,2.91031,2.90691,2.90365,2.90082,2.89822,2.89574,2.89335,2.891,2.88868,2.88632,2.8839,2.88138,2.87871,2.87558,2.87211,2.86857,2.86505,2.86162,2.85868,2.85605,2.85354,2.85112,2.84877,2.84624,2.84362,2.84107,2.8386,2.83624,2.83448,2.83319,2.83185,2.83031,2.82841,2.82571,2.82138,2.81676,2.81205,2.80743,2.80375,2.80093,2.79841,2.79611,2.79393,2.79164,2.78915,2.78666,2.78416,2.78167,2.77917,2.77665,2.77414,2.77163,2.76912,2.76661,2.76411,2.76162,2.75913,2.75664,2.75412,2.7515,2.74891,2.7464,2.74399,2.74176,2.74025,2.7388,2.73731,2.73567,2.73378,2.73067,2.72707,2.72344,2.71993,2.71672,2.71527,2.71438,2.71373,2.71317,2.71253,2.71117,2.70873,2.70614,2.70353,2.70101,2.69902,2.69812,2.69741,2.69676,2.69604,2.69513,2.69339,2.69121,2.68876,2.68606,2.68314,2.67981,2.67626,2.67271,2.66927,2.66603,2.66379,2.66204,2.66047,2.65899,2.65749,2.65557,2.65321,2.65074,2.64818,2.64557,2.64294,2.64032,2.63775,2.63525,2.63287,2.63076,2.62911,2.62754,2.62599,2.62441,2.62271,2.62029,2.61777,2.61521,2.61268,2.61024,2.60847,2.60687,2.60533,2.60377,2.60212,2.6,2.59751,2.59496,2.59241,2.58992,2.58785,2.58622,2.58466,2.58311,2.58151,2.57967,2.57711,2.57449,2.57191,2.56946,2.5673,2.56621,2.56536,2.56465,2.56401,2.56334,2.56233,2.56099,2.5595,2.55784,2.55602,2.55396,2.55151,2.54897,2.54641,2.5439,2.54154,2.53972,2.53803,2.53645,2.53494,2.53346,2.53178,2.53008,2.52842,2.52685,2.52538,2.52425,2.52343,2.52269,2.52196,2.52119,2.52033,2.51894,2.51742,2.5158,2.51412,2.5124,2.51074,2.50912,2.5075,2.50588,2.50426,2.50265,2.50105,2.49945,2.49786,2.49626,2.49466,2.49304,2.49142,2.4898,2.48818,2.48656,2.48496,2.48336,2.48176,2.48016,2.47856,2.47696,2.47534,2.47372,2.4721,2.47048,2.46885,2.46701,2.46523,2.46356,2.46206,2.46076,2.46034,2.46031,2.4604,2.46049,2.46049,2.46028,2.45902,2.45753,2.45588,2.4541,2.45226,2.45041,2.4486,2.44688,2.44531,2.44393,2.44304,2.44281,2.44276,2.44283,2.44293,2.443,2.4426,2.44193,2.44117,2.44034,2.43946,2.43858,2.43779,2.43699,2.4362,2.4354,2.4346,2.43381,2.43301,2.43221,2.43142,2.43062,2.42983,2.42905,2.42828,2.4275,2.42673,2.42595,2.42516,2.42437,2.42358,2.42278,2.42198,2.42118,2.42027,2.41938,2.41853,2.41777,2.4171,2.41674,2.4167,2.41673,2.41678,2.4168,2.41674,2.41627,2.41558,2.41479,2.41394,2.41304,2.41212,2.4112,2.41032,2.40949,2.40874,2.40809,2.40774,2.40761,2.40757,2.4076,2.40768,2.40779,2.40802,2.40821,2.40831,2.40825,2.40798,2.4073,2.40576,2.40407,2.40234,2.40066,2.39914,2.39859,2.39837,2.39834,2.39847,2.39868,2.3989,2.39886,2.39883,2.3988,2.39876,2.39872,2.39869,2.39865,2.39862,2.39858,2.39855,2.39851,2.39848,2.39844,2.3984,2.39837,2.39833,2.3983,2.39828,2.39827,2.39825,2.39823,2.39822,2.3982,2.39817,2.39813,2.3981,2.39806,2.39802,2.39799,2.39795,2.39792,2.39788,2.39785,2.39781,2.39778,2.39774,2.3977,2.39767,2.39763,2.3976,2.39758,2.39757,2.39755,2.39753,2.39752,2.39749,2.39746,2.39743,2.3974,2.39736,2.39732,2.39729,2.39725,2.39722,2.39718,2.39715,2.39711,2.39707,2.39704,2.397,2.39697,2.39693,2.3969,2.39688,2.39687,2.39685,2.39683,2.39682,2.39678,2.39664,2.39652,2.39644,2.39643,2.39651,2.39684,2.39748,2.39818,2.39891,2.39962,2.40028,2.40062,2.40061,2.40054,2.40045,2.40038,2.40038,2.40083,2.4015,2.40221,2.40294,2.40364,2.40427,2.40453,2.4046,2.4046,2.40453,2.40443,2.4043,2.40427,2.40424,2.4042,2.40416,2.40413,2.40406,2.40392,2.4038,2.40373,2.40373,2.40382,2.40419,2.40484,2.40555,2.40628,2.40699,2.40763,2.40792,2.4079,2.40783,2.40774,2.40768,2.40768,2.40817,2.40884,2.40956,2.4103,2.411,2.41162,2.41184,2.41191,2.4119,2.41183,2.41172,2.41158,2.41144,2.41132,2.41125,2.41123,2.4113,2.41161,2.41224,2.41294,2.41367,2.41439,2.41504,2.41547,2.41556,2.41556,2.4155,2.41539,2.41525,2.41519,2.41517,2.41515,2.41514,2.41512,2.4151,2.41497,2.41485,2.41476,2.41473,2.41477,2.41497,2.41559,2.41629,2.41703,2.41775,2.41843,2.41894,2.41906,2.41908,2.41902,2.41892,2.41878,2.41868,2.41865,2.41861,2.41857,2.41854,2.41851,2.41841,2.41829,2.41821,2.41819,2.41824,2.41839,2.41898,2.41966,2.42038,2.42111,2.42179,2.42239,2.42254,2.42258,2.42254,2.42244,2.42231,2.42219,2.42216,2.42212,2.42209,2.42205,2.42202,2.42198,2.42194,2.42191,2.42187,2.42184,2.42181,2.42188,2.42197,2.42203,2.42201,2.42191,2.42168,2.42096,2.42014,2.41929,2.41845,2.41766,2.41717,2.41699,2.41692,2.41692,2.41698,2.41707,2.41709,2.41707,2.41705,2.41704,2.41702,2.417,2.41697,2.41694,2.4169,2.41687,2.41683,2.41679,2.41676,2.41672,2.41669,2.41665,2.41662,2.41658,2.41655,2.41651,2.41648,2.41644,2.41641,2.41647,2.41654,2.41658,2.41655,2.41644,2.41621,2.4155,2.41469,2.41385,2.41302,2.41225,2.41177,2.4116,2.41153,2.41153,2.41159,2.41168,2.41167,2.41163,2.4116,2.41156,2.41153,2.4115,2.41161,2.41169,2.41173,2.4117,2.41158,2.41124,2.41049,2.40966,2.40881,2.40797,2.40721,2.40682,2.40667,2.40662,2.40664,2.4067,2.40679,2.40676,2.40673,2.40669,2.40666,2.40662,2.4066,2.40658,2.40656,2.40654,2.40653,2.40651,2.40649,2.40646,2.40642,2.40639,2.40635,2.40631,2.40636,2.40644,2.40647,2.40644,2.40633,2.4061,2.40539,2.4046,2.40377,2.40294,2.40218,2.40168,2.40151,2.40143,2.40143,2.40149,2.40157,2.40167,2.40174,2.40178,2.40176,2.40164,2.40141,2.4007,2.39989,2.39904,2.3982,2.39741,2.39689,2.39673,2.39667,2.39669,2.39676,2.39686,2.39688,2.39685,2.39681,2.39678,2.39674,2.3967,2.39667,2.39663,2.3966,2.39656,2.39653,2.39651,2.3966,2.39667,2.39668,2.39661,2.39645,2.39602,2.39526,2.39443,2.39359,2.39278,2.39205,2.39178,2.39166,2.39162,2.39165,2.39172,2.39182,2.3919,2.39196,2.39197,2.39191,2.39175,2.39131,2.39056,2.38974,2.38891,2.3881,2.38738,2.38709,2.38696,2.38692,2.38695,2.38702,2.3871,2.38706,2.38703,2.38699,2.38696,2.38692,2.38694,2.38702,2.38707,2.38707,2.38698,2.3868,2.38634,2.38568,2.38492,2.38409,2.38322,2.38232,2.38141,2.38052,2.37968,2.37892,2.37826,2.37785,2.37769,2.37762,2.37763,2.37769,2.37779,2.37802,2.37823,2.37835,2.37833,2.37811,2.37755,2.37604,2.37436,2.37262,2.37093,2.36939,2.36871,2.36845,2.36838,2.36847,2.36867,2.3689,2.36901,2.3691,2.36913,2.3691,2.36897,2.3686,2.36785,2.36702,2.36616,2.36533,2.36457,2.36393,2.36346,2.3632,2.36321,2.36352,2.3642  ;
idx_rfr_Vol73_img = 0.017013,0.018438,0.019129,0.022541,0.027046,0.027542,0.027738,0.029433,0.032607,0.034432,0.034717,0.034863,0.034814,0.034415,0.034118,0.033743,0.033044,0.032163,0.029886,0.026572,0.023714,0.022342,0.022895,0.029880,0.021655,0.016871,0.016988,0.016101,0.015513,0.014854,0.014766,0.014771,0.014618,0.014386,0.014275,0.014029,0.013873,0.013794,0.013616,0.013436,0.013409,0.013316,0.013240,0.013096,0.012844,0.012617,0.012276,0.012017,0.011884,0.011805,0.011739,0.011608,0.011451,0.011160,0.010982,0.010837,0.010608,0.010430,0.010193,0.009949,0.009524,0.009204,0.008906,0.008288,0.008259,0.006893,0.006256,0.004783,0.004980,0.005012,0.004471,0.004473,0.004363,0.004307,0.004309,0.004286,0.004266,0.004305,0.004276,0.004286,0.004292,0.004302,0.004307,0.004353,0.004397,0.004443,0.004489,0.004533,0.004602,0.004669,0.004716,0.004774,0.004948,0.005082,0.005083,0.005270,0.005527,0.005679,0.005762,0.005817,0.005932,0.006055,0.006177,0.006333,0.006691,0.006928,0.007300,0.007507,0.007690,0.007759,0.007936,0.008439,0.008894,0.009233,0.009910,0.010280,0.010576,0.010876,0.011198,0.011673,0.012185,0.013203,0.013453,0.013654,0.013894,0.014060,0.014352,0.014641,0.015030,0.015506,0.015836,0.016224,0.016995,0.017693,0.017935,0.018441,0.018607,0.018989,0.019333,0.019691,0.020120,0.020762,0.021289,0.021843,0.023114,0.023852,0.024423,0.024928,0.025361,0.025618,0.026096,0.026440,0.027160,0.028022,0.028636,0.029519,0.030561,0.031870,0.032667,0.033312,0.033631,0.034173,0.034394,0.034990,0.035713,0.036451,0.037205,0.037973,0.038714,0.039049,0.040462,0.040711,0.041353,0.042553,0.042966,0.043432,0.043547,0.043937,0.044305,0.044254,0.044529,0.044998,0.045798,0.046084,0.046572,0.046858,0.047764,0.048611,0.049900,0.049745,0.050592,0.050617,0.050792,0.051066,0.051051,0.050581,0.050608,0.050407,0.049050,0.048795,0.047173,0.046188,0.045018,0.044007,0.043066,0.042106,0.041865,0.041876,0.042710,0.045052,0.046888,0.047116,0.048958,0.051981,0.056055,0.061754,0.066753,0.069496,0.071746,0.071110,0.057902,0.094201,0.086592,0.088522,0.092026,0.094634,0.100149,0.102806,0.103776,0.104558,0.104971,0.106149,0.10629,0.106267,0.106307,0.105574,0.105314,0.105199,0.103678,0.101258,0.101659,0.100856,0.100148,0.099129,0.097617,0.095271,0.091714,0.090449,0.088781,0.086347,0.085810,0.084481,0.082192,0.080417,0.078370,0.076275,0.075358,0.072422,0.071028,0.068546,0.066224,0.065525,0.064791,0.064560,0.063990,0.063411,0.063429,0.063418,0.063407,0.063470,0.064176,0.064457,0.064910,0.065591,0.066242,0.067249,0.068232,0.068907,0.070235,0.070899,0.072051,0.073028,0.073793,0.075334,0.076890,0.078561,0.078823,0.081817,0.083181,0.084928,0.085804,0.087266,0.089185,0.092035,0.094448,0.095584,0.098292,0.100674,0.10509,0.1076,0.108568,0.110659,0.114265,0.122015,0.125828,0.131309,0.135701,0.13929,0.141691,0.146168,0.151962,0.155577,0.163761,0.171838,0.175816,0.177372,0.180874,0.185595,0.191849,0.195619,0.199675,0.205241,0.222609,0.233777,0.244524,0.252867,0.253985,0.264424,0.277892,0.306018,0.320842,0.326846,0.337086,0.346595,0.351276,0.360086,0.371105,0.376641,0.396459,0.412026,0.423363,0.428527,0.432777,0.439112,0.448633,0.454073,0.459236,0.46889,0.478584,0.488491,0.498568,0.509078,0.517714,0.522484,0.532361,0.533428,0.538829,0.547573,0.551012,0.560564,0.561352,0.567685,0.5695,0.578564,0.589515,0.592256,0.605154,0.617649,0.630448,0.636939,0.64347,0.649762,0.661997,0.664067,0.674279,0.679787,0.695166,0.697174,0.710568,0.717247,0.729089,0.737945,0.772807,0.784678,0.791219,0.797860,0.804065,0.813336,0.831251,0.839201,0.844646,0.853808,0.871996,0.886437,0.894222,0.918693,0.929136,0.939144,0.943991,0.943391,0.942237,0.92733,0.913961,0.896719,0.887175,0.868527,0.845313,0.824644,0.80013,0.789922,0.772608,0.7567,0.740758,0.733402,0.721708,0.705693,0.691852,0.680581,0.661703,0.6477,0.633351,0.600296,0.5757,0.5642,0.552278,0.542367,0.53701,0.526689,0.519232,0.508355,0.502544,0.491719,0.481946,0.475394,0.465349,0.447007,0.440962,0.426193,0.41821,0.413736,0.406762,0.405737,0.395369,0.392975,0.384495,0.379883,0.375216,0.366727,0.36101,0.354893,0.343715,0.339451,0.329435,0.322122,0.320028,0.314479,0.313046,0.309062,0.304971,0.303606,0.297802,0.294736,0.291565,0.288535,0.28249,0.273923,0.26543,0.264521,0.257195,0.254617,0.252103,0.2471,0.247215,0.246222,0.243504,0.238833,0.233619,0.228668,0.223611,0.222896,0.218989,0.217258,0.215354,0.211702,0.211307,0.208915,0.206749,0.204446,0.203813,0.200052,0.197786,0.199024,0.197182,0.194922,0.193936,0.193982,0.193956,0.19375,0.195889,0.195949,0.195478,0.195441,0.19541,0.195377,0.19534,0.195221,0.190544,0.187003,0.183924,0.1807,0.180134,0.178186,0.174872,0.171619,0.170314,0.168583,0.168692,0.168249,0.165744,0.163901,0.162963,0.160134,0.159158,0.156457,0.154955,0.15197,0.15214,0.151291,0.149654,0.146873,0.146062,0.14359,0.142082,0.14057,0.13946,0.138755,0.138206,0.1382,0.136945,0.136851,0.138672,0.140443,0.141836,0.143788,0.146102,0.147522,0.149029,0.148842,0.150148,0.153562,0.154028,0.156965,0.158434,0.160989,0.163133,0.166257,0.167807,0.171066,0.174456,0.176041,0.181461,0.186145,0.187854,0.189781,0.191716,0.193703,0.195783,0.19768,0.201447,0.201534,0.202078,0.204366,0.204895,0.206831,0.208487,0.208232,0.209549,0.211796,0.211814,0.211776,0.21174,0.211829,0.207919,0.208277,0.205705,0.20441,0.204447,0.204505,0.203461,0.201119,0.200859,0.200821,0.201001,0.198124,0.197339,0.197302,0.197381,0.195976,0.195523,0.195443,0.19613,0.197189,0.197105,0.19531,0.19533,0.195291,0.195196,0.196928,0.19679,0.197544,0.19985,0.200143,0.200047,0.200683,0.202966,0.203453,0.203357,0.20388,0.206187,0.206843,0.206961,0.210414,0.210225,0.210188,0.21012,0.211939,0.212661,0.213741,0.213614,0.213577,0.213539,0.213502,0.213466,0.213429,0.213391,0.213354,0.213216,0.21505,0.215074,0.214928,0.216375,0.21516,0.215215,0.216835,0.216682,0.216645,0.216609,0.21657,0.216534,0.216399,0.218278,0.218198,0.219127,0.220155,0.220033,0.219995,0.219947,0.219911,0.219875,0.219836,0.2198,0.219763,0.219727,0.219707,0.219159,0.217771,0.216284,0.215839,0.215741,0.216557,0.217546,0.21924,0.221253,0.221857,0.223151,0.223006,0.222967,0.22292,0.222885,0.222846,0.22281,0.222704,0.223296,0.222643,0.222574,0.224557,0.224346,0.226341,0.226067,0.22829,0.230197,0.230072,0.231437,0.231635,0.234027,0.233746,0.236042,0.237874,0.237692,0.237647,0.237608,0.23757,0.237398,0.239075,0.239475,0.241573,0.241435,0.2414,0.241253,0.245604,0.245415,0.245241,0.247061,0.249642,0.252293,0.253826,0.253548,0.255771,0.255732,0.255554,0.257097,0.257805,0.257982,0.26083,0.2622,0.262028,0.262109,0.264953,0.26638,0.268053,0.268556,0.270461,0.267396,0.290604,0.290604,0.302114,0.302921,0.303762,0.30466,0.305635,0.30671,0.308051,0.309724,0.311495,0.313334,0.315211,0.317096,0.318959,0.320551,0.322033,0.323478,0.324895,0.326293,0.327684,0.329103,0.330574,0.332052,0.333537,0.335027,0.336522,0.338023,0.339601,0.34117,0.342719,0.344236,0.345709,0.347126,0.348331,0.349386,0.350411,0.35143,0.352469,0.353552,0.354773,0.356175,0.357661,0.359228,0.360877,0.362607,0.364431,0.36656,0.368732,0.370913,0.373067,0.375157,0.377149,0.378705,0.379751,0.380752,0.381778,0.382894,0.384168,0.385897,0.388629,0.391601,0.39475,0.398014,0.401331,0.40464,0.407803,0.410298,0.412702,0.415032,0.417309,0.41955,0.421774,0.424025,0.426318,0.428641,0.431006,0.433425,0.43591,0.438473,0.441273,0.444183,0.447166,0.450211,0.453308,0.456446,0.459612,0.462714,0.465834,0.468974,0.472134,0.475313,0.478512,0.481732,0.484977,0.488242,0.491526,0.494828,0.498148,0.501486,0.504836,0.508194,0.511569,0.514964,0.518381,0.52182,0.525282,0.528776,0.532303,0.535856,0.539433,0.543034,0.54666,0.550308,0.554043,0.557842,0.56164,0.565422,0.569174,0.572878,0.576522,0.579781,0.582868,0.585951,0.589074,0.59228,0.595612,0.599177,0.603669,0.608323,0.613083,0.617892,0.622691,0.627424,0.632033,0.635713,0.639235,0.642678,0.646087,0.649508,0.652984,0.656758,0.661055,0.665443,0.66989,0.674359,0.678819,0.683234,0.687267,0.690901,0.69452,0.698175,0.701915,0.705791,0.709854,0.715085,0.720672,0.726362,0.732065,0.737691,0.743153,0.748359,0.752328,0.755679,0.758831,0.76186,0.764842,0.767852,0.771296,0.775588,0.779951,0.784315,0.788607,0.792755,0.796688,0.799789,0.802379,0.80476,0.806978,0.809081,0.811118,0.813531,0.816236,0.81884,0.821278,0.823482,0.825384,0.826635,0.827013,0.827095,0.82695,0.826644,0.826247,0.826398,0.826784,0.827014,0.826994,0.826632,0.825834,0.823231,0.820269,0.817187,0.814173,0.811414,0.810308,0.810028,0.810045,0.810223,0.810421,0.810447,0.809372,0.808108,0.806699,0.805189,0.80362,0.802039,0.800489,0.799007,0.797635,0.796416,0.795415,0.794857,0.79453,0.794428,0.794547,0.794882,0.7955,0.796417,0.797496,0.798701,0.799997,0.801349,0.802723,0.804084,0.805392,0.806612,0.807706,0.80864,0.808934,0.808745,0.808515,0.808349,0.808351,0.808623,0.810127,0.812115,0.814391,0.81689,0.819544,0.822287,0.824613,0.826802,0.829044,0.831367,0.8338,0.836372,0.839311,0.842588,0.846008,0.849546,0.853175,0.856867,0.860549,0.863939,0.867372,0.870875,0.874475,0.878196,0.882065,0.8865,0.891238,0.896075,0.900961,0.905844,0.910675,0.915353,0.919418,0.923365,0.927219,0.931004,0.934744,0.938462,0.942157,0.945873,0.94965,0.953516,0.957501,0.961634,0.966224,0.971544,0.976954,0.982364,0.987684,0.992834,0.997704,1.001244,1.004074,1.006764,1.009424,1.012174,1.015134,1.019294,1.024644,1.030234,1.035944,1.041644,1.047194,1.052484,1.056524,1.060064,1.063264,1.066154,1.068744,1.071064,1.073044,1.074794,1.076374,1.077824,1.079184,1.080494,1.082214,1.083984,1.085674,1.087234,1.088614,1.089774,1.090464,1.090844,1.090934,1.090724,1.090204,1.089324,1.087854,1.086144,1.084234,1.082204,1.080104,1.078434,1.076884,1.075234,1.073414,1.071364,1.068724,1.064914,1.060994,1.057164,1.053594,1.050464,1.050014,1.050034,1.050264,1.050464,1.050384,1.049174,1.045904,1.042254,1.038394,1.034524,1.030924,1.028724,1.026814,1.025134,1.023604,1.022174,1.020764,1.019314,1.017774,1.016064,1.014144,1.011814,1.008424,1.004844,1.001214,0.997644,0.994274,0.992034,0.990154,0.988494,0.986994,0.985584,0.984204,0.982784,0.981284,0.979634,0.977794,0.975664,0.972224,0.968644,0.965104,0.961754,0.958781,0.957799,0.957748,0.957938,0.958146,0.958152,0.957635,0.955004,0.951916,0.948484,0.944823,0.941047,0.937493,0.934042,0.93071,0.927552,0.924624,0.9223,0.920475,0.918874,0.917437,0.916107,0.914825,0.913516,0.912146,0.910661,0.909006,0.907128,0.904299,0.900989,0.89766,0.894466,0.891565,0.889891,0.889726,0.889853,0.890066,0.890157,0.889919,0.887866,0.884916,0.881708,0.878398,0.875145,0.872638,0.87088,0.869345,0.867976,0.866719,0.865515,0.864299,0.863029,0.861652,0.860115,0.858365,0.855807,0.852649,0.849457,0.84638,0.843571,0.84171,0.841259,0.841173,0.84131,0.841524,0.841673,0.840974,0.839735,0.838327,0.836797,0.835188,0.833588,0.83217,0.830755,0.829341,0.827928,0.826516,0.825098,0.823679,0.822261,0.820845,0.819433,0.817966,0.81637,0.814833,0.813396,0.812102,0.810995,0.810848,0.811021,0.8112,0.811249,0.811032,0.810246,0.807614,0.804708,0.801706,0.798792,0.796144,0.795078,0.794657,0.794584,0.794769,0.795121,0.795476,0.795424,0.795372,0.795319,0.795266,0.795213,0.79526,0.795409,0.795497,0.795481,0.795322,0.794976,0.79406,0.792864,0.791513,0.790051,0.78852,0.786965,0.785431,0.783954,0.782575,0.781335,0.780276,0.779794,0.779576,0.779515,0.779571,0.779703,0.779836,0.779785,0.779735,0.779684,0.779633,0.779582,0.779531,0.77948,0.77943,0.779379,0.779328,0.779277,0.779224,0.779172,0.779119,0.779066,0.779014,0.778961,0.77891,0.778859,0.778808,0.778757,0.778706,0.778656,0.778605,0.778554,0.778503,0.778452,0.778401,0.77835,0.7783,0.778249,0.778198,0.778147,0.778096,0.778045,0.777994,0.777943,0.777892,0.777841,0.777791,0.77774,0.777689,0.777639,0.777588,0.777536,0.777484,0.777432,0.777379,0.777326,0.777273,0.777221,0.777169,0.777118,0.777067,0.777017,0.776966,0.776915,0.776865,0.776814,0.776763,0.776712,0.776661,0.77661,0.776559,0.776508,0.776457,0.776406,0.776356,0.776305,0.776254,0.776203,0.776152,0.776101,0.77605,0.775999,0.775948,0.775898,0.775847,0.775796,0.775745,0.775694,0.775643,0.775592,0.775541,0.77549,0.77544,0.775389,0.775338,0.775287,0.775236,0.775185,0.775134,0.775083,0.775032,0.774981,0.774931,0.77488,0.774829,0.774778,0.774727,0.774676,0.774625,0.774574,0.774523,0.774473,0.774422,0.774371,0.77432,0.774269,0.774218,0.774167,0.774116,0.774065,0.774014,0.773964,0.773913,0.773862,0.773811,0.77376,0.773817,0.773966,0.774055,0.774041,0.773884,0.773543,0.772488,0.771143,0.769722,0.768307,0.766981,0.766058,0.765748,0.765616,0.765621,0.765721,0.765877,0.765901,0.765852,0.765803,0.765754,0.765705,0.765655,0.765808,0.765929,0.76597,0.765893,0.765658,0.765056,0.763809,0.762445,0.761043,0.759684,0.758448,0.758066,0.758023,0.758066,0.758115,0.758089,0.75783,0.756624,0.755288,0.753901,0.752542,0.75129,0.750729,0.750663,0.750696,0.750749,0.750742,0.750595,0.749678,0.748529,0.747239,0.745847,0.744393,0.743001,0.741714,0.740429,0.739145,0.737864,0.73659,0.735543,0.734455,0.73328,0.731971,0.730481,0.728327,0.725624,0.722886,0.720244,0.717826,0.716171,0.715771,0.715687,0.715799,0.715982,0.716113,0.71555,0.714494,0.713292,0.711984,0.710607,0.709228,0.70801,0.706795,0.705581,0.704369,0.703159,0.701952,0.700748,0.699545,0.698343,0.697142,0.695904,0.694525,0.693192,0.691941,0.690812,0.689841,0.689671,0.689813,0.689967,0.690016,0.689844,0.689236,0.686993,0.684508,0.681937,0.679435,0.677155,0.676336,0.676121,0.676145,0.676293,0.67645,0.676412,0.675499,0.67443,0.673241,0.671966,0.670643,0.669305,0.66799,0.666734,0.665575,0.664547,0.663768,0.66347,0.663334,0.663323,0.6634,0.663531,0.663787,0.664106,0.664312,0.66433,0.664086,0.663505,0.661633,0.659281,0.656807,0.65436,0.65209,0.650765,0.650316,0.650178,0.650274,0.65053,0.650872,0.651046,0.651158,0.651207,0.651156,0.65097,0.650558,0.649655,0.648602,0.647434,0.646188,0.6449,0.643614,0.642359,0.641166,0.640069,0.639101,0.638432,0.638328,0.638333,0.63838,0.638401,0.638326,0.6377,0.636615,0.635451,0.634274,0.633153,0.632207,0.632077,0.632067,0.632111,0.632141,0.632088,0.631622,0.630569,0.629426,0.628258,0.627133,0.626117,0.625735,0.625564,0.625519,0.625568,0.625676,0.625744,0.625556,0.625403,0.625313,0.625315,0.625439,0.626161,0.627434,0.628686,0.629787,0.630604,0.631008,0.629978,0.627874,0.625519,0.623083,0.620742,0.619128,0.618634,0.618452,0.618512,0.618739,0.619063,0.619146,0.619106,0.619066,0.619025,0.618985,0.618945,0.618903,0.618861,0.618818,0.618776,0.618734,0.618692,0.618652,0.618612,0.618571,0.618531,0.618491,0.618449,0.618407,0.618365,0.618323,0.618281,0.618239,0.618198,0.618158,0.618117,0.618077,0.618037,0.617996,0.617954,0.617912,0.61787,0.617827,0.617785,0.61783,0.617948,0.618018,0.618007,0.617882,0.617611,0.616766,0.615692,0.614555,0.613422,0.612358,0.611589,0.611336,0.611225,0.611224,0.611301,0.611423,0.611448,0.611406,0.611364,0.611322,0.611279,0.611237,0.611196,0.611156,0.611116,0.611075,0.611035,0.610995,0.610955,0.610914,0.610874,0.610834,0.610793,0.610753,0.610713,0.610672,0.610632,0.610591,0.610551,0.610511,0.610471,0.610431,0.61039,0.61035,0.610309,0.610267,0.610225,0.610182,0.61014,0.610098,0.610056,0.610016,0.609975,0.609935,0.609895,0.609855,0.609815,0.609774,0.609734,0.609693,0.609653,0.609613,0.609572,0.609532,0.609492,0.609451,0.609411,0.609371,0.60933,0.60929,0.609249,0.609209,0.609169,0.609128,0.609088,0.609048,0.609007,0.608967,0.608927,0.608886,0.608846,0.608806,0.608766,0.608725,0.608648,0.608462,0.608312,0.608224,0.608227,0.60835,0.608876,0.609755,0.610713,0.611695,0.612645,0.613505,0.613929,0.614032,0.61402,0.613922,0.613765,0.613578,0.613527,0.613487,0.613447,0.613406,0.613366,0.613324,0.613282,0.61324,0.613198,0.613156,0.613114,0.613072,0.613032,0.612991,0.612951,0.612911,0.612871,0.612831,0.612791,0.61275,0.61271,0.612669,0.612628,0.612586,0.612544,0.612502,0.61246,0.612418,0.612376,0.612336,0.612295,0.612255,0.612215,0.612175,0.612134,0.612094,0.612054,0.612013,0.611973,0.611927,0.611739,0.61158,0.611479,0.611464,0.611563,0.611965,0.612824,0.613775,0.61476,0.615724,0.61661,0.617162,0.617292,0.617302,0.617219,0.617071,0.616887,0.616804,0.616762,0.616719,0.616677,0.616635,0.616593,0.616552,0.616512,0.616471,0.616431,0.616391,0.616351,0.616311,0.616271,0.61623,0.61619,0.616149,0.616012,0.615835,0.615705,0.615649,0.615697,0.615876,0.616655,0.617582,0.618567,0.619554,0.620485,0.621298,0.621485,0.621539,0.621488,0.621361,0.621186,0.620993,0.620811,0.620665,0.620585,0.620599,0.620734,0.621313,0.622208,0.623179,0.624171,0.625127,0.625991,0.626402,0.6265,0.626485,0.626383,0.626224,0.626034,0.62584,0.625673,0.625562,0.625537,0.625625,0.626296,0.628378,0.630291,0.631752,0.632475,0.632175,0.629457,0.623422,0.616874,0.610292,0.604154,0.60124,0.600076,0.599848,0.600361,0.601421,0.602754,0.603415,0.604209,0.605109,0.606088,0.607118,0.608053,0.608427,0.608913,0.609604,0.610596,0.611982,0.614408,0.61904,0.624085,0.629327,0.63455,0.639536,0.64407,0.647643,0.648515,0.648829,0.648707,0.64827,0.647641,0.647225,0.647181,0.647137,0.647093,0.647049,0.647006,0.646963,0.646921,0.646879,0.646837,0.646795,0.646753,0.646709,0.646665,0.646621,0.646577,0.646533,0.64649,0.646447,0.646405,0.646363,0.646321,0.646279,0.646136,0.645954,0.64582,0.645764,0.645817,0.646007,0.646826,0.647795,0.648824,0.649854,0.650826,0.651666,0.651705,0.651636,0.65152,0.651415,0.651379,0.651688,0.652598,0.653606,0.654652,0.655676,0.656618,0.657214,0.657354,0.657364,0.657276,0.65712,0.656924,0.656833,0.656789,0.656745,0.656701,0.656657,0.656612,0.65641,0.656238,0.656127,0.656107,0.656208,0.656565,0.657316,0.658205,0.659202,0.660278,0.661402,0.662547,0.663684,0.664781,0.665806,0.66673,0.667522,0.667991,0.668123,0.668127,0.668032,0.66787,0.66767,0.66759,0.667546,0.667502,0.667458,0.667414,0.66737,0.667327,0.667283,0.667239,0.667196,0.667151,0.66699,0.666663,0.666413,0.666299,0.666376,0.666701,0.668012,0.669909,0.671967,0.674071,0.676109,0.677967,0.679709,0.681191,0.68205,0.682111,0.681198;
}

// $Id$
// ncgen -b -o ${DATA}/aca/idx_rfr_triaud_Fe2O3.nc ${HOME}/idx_rfr/idx_rfr_triaud_Fe2O3.cdl

netcdf idx_rfr_triaud_Fe2O3 {
dimensions:
	bnd = UNLIMITED ; // (801 currently)
variables:

// global attributes:
	:history = "Thu Jan 26 22:19:38 2006: ncrename -O -d u,bnd idx_rfr_triaud_Fe2O3.nc" ;
	:source="
Database of Optical Constants for Cosmic Dust (DOCCD)
Laboratory Astrophysics Group of the AIU Jena 
http://www.astro.uni-jena.de/Laboratory/OCDB/oxsul.html
Iron oxides, created by Amaury Triaud <at42@st-andrews.ac.uk> unpublished
Charlie Zender <zender@uci.edu> standardized 20060129.

As mentioned at web-site, these data appear to be E-ray (rather than O-ray)
Measurements by Shettle have both E-ray and O-ray

Procedure to create netCDF from text file:
fl_txt=idx_rfr_triaud_Fe2O3
cat > /tmp/${fl_txt}.header << EOF
bnd:f idx_rfr_Fe2O3_rl:f idx_rfr_Fe2O3_img:f
EOF
tbl2cdf -h /tmp/${fl_txt}.header ~/idx_rfr/doccd/idx_rfr_fe2o3.txt ~/idx_rfr/${fl_txt}.nc
ncrename -O -d u,bnd ${fl_txt}.nc
ncks ~/idx_rfr/${fl_txt}.nc | m
ncdump ~/idx_rfr/${fl_txt}.nc > ~/idx_rfr/${fl_txt}.cdl
";

	float bnd(bnd);
	bnd:long_name = "Band center wavelength";
	bnd:units = "micron";
	bnd:C_format = "%.5g";

	float idx_rfr_Fe2O3_doccd_rl(bnd);
	idx_rfr_Fe2O3_doccd_rl:long_name = "Hematite real index of refraction E-ray";
	idx_rfr_Fe2O3_doccd_rl:units = "";
	idx_rfr_Fe2O3_doccd_rl:composition = "Fe2O3";
	idx_rfr_Fe2O3_doccd_rl:C_format = "%.4g";

	float idx_rfr_Fe2O3_doccd_img(bnd);
	idx_rfr_Fe2O3_doccd_img:long_name = "Hematite imaginary index of refraction E-ray";
	idx_rfr_Fe2O3_doccd_img:units = "";
	idx_rfr_Fe2O3_doccd_img:composition = "Fe2O3";
	idx_rfr_Fe2O3_doccd_img:C_format = "%.3g";

data:

 bnd = 0.1, 0.10116, 0.10233, 0.10351, 0.10471, 0.10593, 0.10715, 0.10839, 
    0.10965, 0.11092, 0.1122, 0.1135, 0.11482, 0.11614, 0.11749, 0.11885, 
    0.12023, 0.12162, 0.12303, 0.12445, 0.12589, 0.12735, 0.12882, 0.13032, 
    0.13183, 0.13335, 0.1349, 0.13646, 0.13804, 0.13964, 0.14125, 0.14289, 
    0.14454, 0.14622, 0.14791, 0.14962, 0.15136, 0.15311, 0.15488, 0.15668, 
    0.15849, 0.16032, 0.16218, 0.16406, 0.16596, 0.16788, 0.16982, 0.17179, 
    0.17378, 0.17579, 0.17783, 0.17989, 0.18197, 0.18408, 0.18621, 0.18836, 
    0.19055, 0.19275, 0.19498, 0.19724, 0.19953, 0.20184, 0.20417, 0.20654, 
    0.20893, 0.21135, 0.2138, 0.21627, 0.21878, 0.22131, 0.22387, 0.22646, 
    0.22909, 0.23174, 0.23442, 0.23714, 0.23988, 0.24266, 0.24547, 0.24831, 
    0.25119, 0.2541, 0.25704, 0.26002, 0.26303, 0.26607, 0.26915, 0.27227, 
    0.27542, 0.27861, 0.28184, 0.2851, 0.2884, 0.29174, 0.29512, 0.29854, 
    0.302, 0.30549, 0.30903, 0.31261, 0.31623, 0.31989, 0.32359, 0.32734, 
    0.33113, 0.33497, 0.33884, 0.34277, 0.34674, 0.35075, 0.35481, 0.35892, 
    0.36308, 0.36728, 0.37154, 0.37584, 0.38019, 0.38459, 0.38905, 0.39355, 
    0.39811, 0.40272, 0.40738, 0.4121, 0.41687, 0.4217, 0.42658, 0.43152, 
    0.43652, 0.44157, 0.44668, 0.45186, 0.45709, 0.46238, 0.46774, 0.47315, 
    0.47863, 0.48417, 0.48978, 0.49545, 0.50119, 0.50699, 0.51286, 0.5188, 
    0.52481, 0.53088, 0.53703, 0.54325, 0.54954, 0.5559, 0.56234, 0.56885, 
    0.57544, 0.5821, 0.58884, 0.59566, 0.60256, 0.60954, 0.6166, 0.62373, 
    0.63096, 0.63826, 0.64565, 0.65313, 0.66069, 0.66834, 0.67608, 0.68391, 
    0.69183, 0.69984, 0.70795, 0.71614, 0.72444, 0.73282, 0.74131, 0.74989, 
    0.75858, 0.76736, 0.77625, 0.78524, 0.79433, 0.80353, 0.81283, 0.82224, 
    0.83176, 0.8414, 0.85114, 0.86099, 0.87096, 0.88105, 0.89125, 0.90157, 
    0.91201, 0.92257, 0.93325, 0.94406, 0.95499, 0.96605, 0.97724, 0.98855, 
    1, 1.01158, 1.02329, 1.03514, 1.04713, 1.05925, 1.07152, 1.08393, 
    1.09648, 1.10917, 1.12202, 1.13501, 1.14815, 1.16145, 1.1749, 1.1885, 
    1.20226, 1.21619, 1.23027, 1.24451, 1.25893, 1.2735, 1.28825, 1.30317, 
    1.31826, 1.33352, 1.34896, 1.36458, 1.38038, 1.39637, 1.41254, 1.42889, 
    1.44544, 1.46218, 1.47911, 1.49624, 1.51356, 1.53109, 1.54882, 1.56675, 
    1.58489, 1.60325, 1.62181, 1.64059, 1.65959, 1.6788, 1.69824, 1.71791, 
    1.7378, 1.75792, 1.77828, 1.79887, 1.8197, 1.84077, 1.86209, 1.88365, 
    1.90546, 1.92752, 1.94984, 1.97242, 1.99526, 2.01837, 2.04174, 2.06538, 
    2.0893, 2.11349, 2.13796, 2.16272, 2.18776, 2.21309, 2.23872, 2.26464, 
    2.29087, 2.31739, 2.34423, 2.37137, 2.39883, 2.42661, 2.45471, 2.48313, 
    2.51189, 2.54097, 2.5704, 2.60016, 2.63027, 2.66073, 2.69153, 2.7227, 
    2.75423, 2.78612, 2.81838, 2.85102, 2.88403, 2.91743, 2.95121, 2.98538, 
    3.01995, 3.05492, 3.0903, 3.12608, 3.16228, 3.1989, 3.23594, 3.27341, 
    3.31131, 3.34965, 3.38844, 3.42768, 3.46737, 3.50752, 3.54813, 3.58922, 
    3.63078, 3.67282, 3.71535, 3.75837, 3.80189, 3.84592, 3.89045, 3.9355, 
    3.98107, 4.02717, 4.0738, 4.12098, 4.16869, 4.21697, 4.2658, 4.31519, 
    4.36516, 4.4157, 4.46684, 4.51856, 4.57088, 4.62381, 4.67735, 4.73151, 
    4.7863, 4.84172, 4.89779, 4.9545, 5.01187, 5.06991, 5.12861, 5.188, 
    5.24807, 5.30884, 5.37032, 5.4325, 5.49541, 5.55904, 5.62341, 5.68853, 
    5.7544, 5.82103, 5.88844, 5.95662, 6.0256, 6.09537, 6.16595, 6.23735, 
    6.30957, 6.38263, 6.45654, 6.53131, 6.60693, 6.68344, 6.76083, 6.83912, 
    6.91831, 6.99842, 7.07946, 7.16143, 7.24436, 7.32825, 7.4131, 7.49894, 
    7.58578, 7.67361, 7.76247, 7.85236, 7.94328, 8.03526, 8.12831, 8.22243, 
    8.31764, 8.41395, 8.51138, 8.60994, 8.70964, 8.81049, 8.91251, 9.01571, 
    9.12011, 9.22571, 9.33254, 9.44061, 9.54993, 9.66051, 9.77237, 9.88553, 
    10, 10.11579, 10.23293, 10.35142, 10.47129, 10.59254, 10.71519, 10.83927, 
    10.96478, 11.09175, 11.22018, 11.35011, 11.48154, 11.61449, 11.74898, 
    11.88502, 12.02264, 12.16186, 12.30269, 12.44515, 12.58925, 12.73503, 
    12.8825, 13.03167, 13.18257, 13.33521, 13.48963, 13.64583, 13.80384, 
    13.96368, 14.12538, 14.28894, 14.4544, 14.62177, 14.79108, 14.96236, 
    15.13561, 15.31087, 15.48817, 15.66751, 15.84893, 16.03245, 16.2181, 
    16.4059, 16.59587, 16.78804, 16.98244, 17.17908, 17.37801, 17.57924, 
    17.78279, 17.98871, 18.19701, 18.40772, 18.62087, 18.83649, 19.05461, 
    19.27525, 19.49845, 19.72423, 19.95262, 20.18366, 20.41738, 20.6538, 
    20.89296, 21.13489, 21.37962, 21.62719, 21.87762, 22.13095, 22.38721, 
    22.64644, 22.90868, 23.17395, 23.44229, 23.71374, 23.98833, 24.2661, 
    24.54709, 24.83133, 25.11886, 25.40973, 25.70396, 26.0016, 26.30268, 
    26.60725, 26.91535, 27.22701, 27.54229, 27.86121, 28.18383, 28.51018, 
    28.84032, 29.17427, 29.51209, 29.85383, 30.19952, 30.54921, 30.90295, 
    31.26079, 31.62278, 31.98895, 32.35937, 32.73407, 33.11311, 33.49654, 
    33.88442, 34.27678, 34.67369, 35.07519, 35.48134, 35.89219, 36.30781, 
    36.72823, 37.15352, 37.58374, 38.01894, 38.45918, 38.90451, 39.35501, 
    39.81072, 40.2717, 40.73803, 41.20975, 41.68694, 42.16965, 42.65795, 
    43.15191, 43.65158, 44.15704, 44.66836, 45.18559, 45.70882, 46.2381, 
    46.77351, 47.31513, 47.86301, 48.41724, 48.97788, 49.54502, 50.11872, 
    50.69907, 51.28614, 51.88, 52.48075, 53.08844, 53.70318, 54.32503, 
    54.95409, 55.59043, 56.23413, 56.88529, 57.54399, 58.21032, 58.88437, 
    59.56621, 60.25596, 60.95369, 61.6595, 62.37348, 63.09573, 63.82635, 
    64.56542, 65.31306, 66.06934, 66.83439, 67.6083, 68.39116, 69.1831, 
    69.9842, 70.79458, 71.61434, 72.4436, 73.28245, 74.13102, 74.98942, 
    75.85776, 76.73615, 77.62471, 78.52356, 79.43282, 80.35261, 81.28305, 
    82.22426, 83.17638, 84.13951, 85.1138, 86.09938, 87.09636, 88.10489, 
    89.12509, 90.15711, 91.20108, 92.25714, 93.32543, 94.40609, 95.49926, 
    96.60509, 97.72372, 98.85531, 100, 101.158, 102.3293, 103.5142, 104.7129, 
    105.9254, 107.1519, 108.3927, 109.6478, 110.9175, 112.2019, 113.5011, 
    114.8154, 116.1449, 117.4898, 118.8502, 120.2264, 121.6186, 123.0269, 
    124.4515, 125.8925, 127.3503, 128.825, 130.3167, 131.8257, 133.3521, 
    134.8963, 136.4583, 138.0384, 139.6368, 141.2538, 142.8894, 144.544, 
    146.2177, 147.9108, 149.6236, 151.3561, 153.1087, 154.8817, 156.6751, 
    158.4893, 160.3245, 162.181, 164.059, 165.9587, 167.8804, 169.8244, 
    171.7908, 173.7801, 175.7924, 177.8279, 179.8871, 181.9701, 184.0772, 
    186.2087, 188.3649, 190.5461, 192.7525, 194.9845, 197.2423, 199.5262, 
    201.8366, 204.1738, 206.538, 208.9296, 211.3489, 213.7962, 216.2719, 
    218.7762, 221.3095, 223.8721, 226.4644, 229.0868, 231.7395, 234.4229, 
    237.1374, 239.8833, 242.661, 245.4709, 248.3133, 251.1886, 254.0973, 
    257.0396, 260.016, 263.0268, 266.0725, 269.1535, 272.2701, 275.4229, 
    278.6121, 281.8383, 285.1018, 288.4031, 291.7427, 295.1209, 298.5383, 
    301.9952, 305.4921, 309.0295, 312.6079, 316.2278, 319.8895, 323.5937, 
    327.3407, 331.1311, 334.9655, 338.8441, 342.7678, 346.7368, 350.7519, 
    354.8134, 358.9219, 363.0781, 367.2823, 371.5352, 375.8374, 380.1894, 
    384.5918, 389.0451, 393.5501, 398.1072, 402.717, 407.3803, 412.0975, 
    416.8694, 421.6965, 426.5795, 431.5191, 436.5158, 441.5705, 446.6836, 
    451.8559, 457.0882, 462.381, 467.7351, 473.1512, 478.6301, 484.1724, 
    489.7788, 495.4502, 501.1872, 506.9907, 512.8614, 518.8, 524.8074, 
    530.8845, 537.0318, 543.2503, 549.5409, 555.9042, 562.3413, 568.8529, 
    575.4399, 582.1032, 588.8437, 595.6622, 602.5596, 609.5369, 616.595, 
    623.7349, 630.9573, 638.2635, 645.6542, 653.1306, 660.6934, 668.3439, 
    676.083, 683.9116, 691.831, 699.842, 707.9458, 716.1434, 724.436, 
    732.8245, 741.3102, 749.8942, 758.5776, 767.3615, 776.2471, 785.2357, 
    794.3282, 803.5261, 812.8305, 822.2427, 831.7638, 841.3951, 851.1381, 
    860.9938, 870.9636, 881.0489, 891.2509, 901.5712, 912.0109, 922.5714, 
    933.2543, 944.0609, 954.9926, 966.0509, 977.2372, 988.5531, 1000 ;

 idx_rfr_Fe2O3_doccd_rl = 1.78002, 1.76602, 1.75226, 1.73873, 1.72539, 1.71223, 
    1.69921, 1.68633, 1.67357, 1.66091, 1.64832, 1.6358, 1.62333, 1.61089, 
    1.5985, 1.58611, 1.57372, 1.56134, 1.54896, 1.53655, 1.52414, 1.51171, 
    1.49927, 1.48682, 1.47437, 1.46195, 1.44955, 1.4372, 1.42494, 1.41278, 
    1.40077, 1.38897, 1.37741, 1.36616, 1.3553, 1.3449, 1.33506, 1.32586, 
    1.31744, 1.30987, 1.3033, 1.29783, 1.2936, 1.29072, 1.2893, 1.28943, 
    1.29122, 1.29474, 1.30003, 1.30713, 1.31606, 1.32682, 1.33936, 1.35366, 
    1.36964, 1.38718, 1.40622, 1.42658, 1.44816, 1.47077, 1.49424, 1.51839, 
    1.54301, 1.56792, 1.5929, 1.61776, 1.64228, 1.66629, 1.68962, 1.71212, 
    1.73365, 1.75411, 1.77342, 1.79155, 1.80848, 1.82425, 1.83892, 1.85259, 
    1.8654, 1.87752, 1.88918, 1.90059, 1.91203, 1.92375, 1.93603, 1.9491, 
    1.96316, 1.97833, 1.99463, 2.01195, 2.03006, 2.04857, 2.06696, 2.08466, 
    2.10101, 2.11541, 2.12726, 2.1361, 2.14161, 2.14397, 2.14532, 2.15664, 
    2.19727, 2.21595, 2.20136, 2.18394, 2.16891, 2.15612, 2.14537, 2.13686, 
    2.13104, 2.12857, 2.13022, 2.13684, 2.14928, 2.16832, 2.19459, 2.22848, 
    2.27003, 2.31884, 2.37399, 2.43408, 2.49723, 2.56126, 2.62382, 2.68272, 
    2.73604, 2.78242, 2.82103, 2.85166, 2.8746, 2.89056, 2.90064, 2.9062, 
    2.90901, 2.91125, 2.91566, 2.92534, 2.94301, 2.9694, 3.00155, 3.03298, 
    3.05697, 3.06997, 3.07238, 3.06671, 3.0558, 3.04192, 3.02662, 3.01086, 
    2.9952, 2.97995, 2.96528, 2.95125, 2.93787, 2.92515, 2.91307, 2.90157, 
    2.89064, 2.88024, 2.87033, 2.86089, 2.85188, 2.84328, 2.83505, 2.82719, 
    2.81966, 2.81243, 2.80552, 2.79888, 2.7925, 2.78637, 2.78048, 2.77481, 
    2.76935, 2.7641, 2.75903, 2.75415, 2.74943, 2.74488, 2.74049, 2.73624, 
    2.73214, 2.72818, 2.72434, 2.72063, 2.71703, 2.71355, 2.71018, 2.70692, 
    2.70375, 2.70068, 2.6977, 2.69482, 2.69201, 2.68929, 2.68664, 2.68408, 
    2.68158, 2.67915, 2.67679, 2.6745, 2.67226, 2.67009, 2.66798, 2.66592, 
    2.66392, 2.66196, 2.66006, 2.65821, 2.6564, 2.65463, 2.65292, 2.65124, 
    2.64961, 2.64801, 2.64644, 2.64492, 2.64343, 2.64197, 2.64055, 2.63916, 
    2.6378, 2.63647, 2.63517, 2.63389, 2.63264, 2.63142, 2.63022, 2.62904, 
    2.62788, 2.62675, 2.62564, 2.62455, 2.62348, 2.62242, 2.62139, 2.62037, 
    2.61937, 2.61838, 2.61742, 2.61646, 2.61552, 2.6146, 2.61367, 2.61277, 
    2.61188, 2.611, 2.61013, 2.60926, 2.60841, 2.60757, 2.60674, 2.60592, 
    2.6051, 2.60428, 2.60348, 2.60268, 2.60187, 2.60108, 2.6003, 2.59951, 
    2.59874, 2.59796, 2.59718, 2.59641, 2.59564, 2.59487, 2.5941, 2.59333, 
    2.59255, 2.59179, 2.59101, 2.59024, 2.58946, 2.58869, 2.5879, 2.58711, 
    2.58633, 2.58553, 2.58473, 2.58393, 2.58312, 2.5823, 2.58148, 2.58065, 
    2.57981, 2.57896, 2.57811, 2.57725, 2.57637, 2.57549, 2.57459, 2.57368, 
    2.57277, 2.57183, 2.57089, 2.56993, 2.56895, 2.56797, 2.56697, 2.56595, 
    2.56492, 2.56387, 2.5628, 2.56171, 2.5606, 2.55948, 2.55834, 2.55717, 
    2.55598, 2.55477, 2.55354, 2.55228, 2.551, 2.54969, 2.54835, 2.54699, 
    2.5456, 2.54418, 2.54273, 2.54125, 2.53974, 2.5382, 2.53662, 2.53501, 
    2.53336, 2.53167, 2.52994, 2.52818, 2.52638, 2.52453, 2.52265, 2.52072, 
    2.51874, 2.51672, 2.51464, 2.51252, 2.51035, 2.50812, 2.50585, 2.50351, 
    2.50111, 2.49866, 2.49614, 2.49357, 2.49092, 2.48821, 2.48544, 2.48259, 
    2.47966, 2.47667, 2.47359, 2.47043, 2.46718, 2.46386, 2.46045, 2.45694, 
    2.45333, 2.44963, 2.44584, 2.44193, 2.43792, 2.4338, 2.42956, 2.42521, 
    2.42073, 2.41612, 2.41138, 2.40651, 2.4015, 2.39635, 2.39103, 2.38557, 
    2.37993, 2.37414, 2.36817, 2.36202, 2.35568, 2.34914, 2.3424, 2.33545, 
    2.32829, 2.32089, 2.31326, 2.30537, 2.29724, 2.28883, 2.28014, 2.27116, 
    2.26187, 2.25227, 2.24234, 2.23204, 2.22139, 2.21035, 2.1989, 2.18704, 
    2.17475, 2.16195, 2.14868, 2.1349, 2.12058, 2.10565, 2.09013, 2.07396, 
    2.05708, 2.03951, 2.02112, 2.00193, 1.98185, 1.96081, 1.93878, 1.91562, 
    1.89134, 1.86574, 1.83879, 1.81037, 1.78026, 1.74852, 1.71463, 1.67869, 
    1.64047, 1.59933, 1.55538, 1.50823, 1.45679, 1.4011, 1.34049, 1.27377, 
    1.1992, 1.1159, 1.02175, 0.9138, 0.78681, 0.63808, 0.4838, 0.36478, 
    0.29768, 0.26348, 0.24605, 0.23804, 0.23632, 0.23968, 0.24741, 0.2597, 
    0.27724, 0.30131, 0.33404, 0.37891, 0.44171, 0.53228, 0.66797, 0.87984, 
    1.23932, 1.83124, 2.56942, 2.99043, 2.91284, 2.50529, 1.99266, 1.51275, 
    1.15238, 0.96852, 0.89396, 0.89879, 0.97789, 1.14105, 1.43073, 2.00875, 
    3.04434, 4.48713, 6.20539, 6.54074, 6.26921, 5.72129, 5.16372, 4.70047, 
    4.2824, 3.90256, 3.5591, 3.22627, 2.89665, 2.56049, 2.20253, 1.83298, 
    1.45146, 1.14984, 0.90227, 0.79439, 0.71816, 0.68068, 0.67364, 0.67778, 
    0.70695, 0.75028, 0.81185, 0.90687, 1.01622, 1.20653, 1.42616, 1.81809, 
    2.35818, 3.2998, 4.86014, 7.42477, 9.77892, 11.8768, 12.60913, 11.84317, 
    11.07721, 10.31125, 9.64452, 9.13392, 8.6659, 8.31298, 7.9691, 7.70796, 
    7.44682, 7.22949, 7.01864, 6.81216, 6.60879, 6.35915, 5.96098, 5.56281, 
    6.17723, 7.00697, 7.41442, 7.01229, 6.61016, 6.42921, 6.30779, 6.19339, 
    6.11706, 6.04074, 5.97292, 5.91589, 5.85885, 5.80916, 5.76362, 5.71809, 
    5.67848, 5.64092, 5.60337, 5.5703, 5.53875, 5.50719, 5.4787, 5.45188, 
    5.42506, 5.39989, 5.37692, 5.35395, 5.33126, 5.31148, 5.2917, 5.27192, 
    5.25378, 5.23669, 5.2196, 5.20251, 5.18768, 5.17287, 5.15807, 5.14368, 
    5.13084, 5.118, 5.10516, 5.09277, 5.08163, 5.07049, 5.05935, 5.04841, 
    5.03875, 5.02909, 5.01943, 5.00978, 5.00114, 4.99278, 4.98442, 4.97606, 
    4.96794, 4.96072, 4.95349, 4.94627, 4.93905, 4.93222, 4.926, 4.91978, 
    4.91356, 4.90734, 4.90137, 4.89604, 4.8907, 4.88537, 4.88004, 4.8747, 
    4.87003, 4.86549, 4.86094, 4.85639, 4.85184, 4.84733, 4.84347, 4.83962, 
    4.83576, 4.8319, 4.82805, 4.82419, 4.82086, 4.81762, 4.81437, 4.81113, 
    4.80789, 4.80465, 4.80149, 4.79879, 4.79609, 4.79339, 4.79069, 4.78799, 
    4.78529, 4.78259, 4.78033, 4.77811, 4.77588, 4.77366, 4.77144, 4.76922, 
    4.76699, 4.76478, 4.76298, 4.76117, 4.75937, 4.75756, 4.75576, 4.75396, 
    4.75215, 4.75035, 4.74866, 4.74723, 4.74579, 4.74436, 4.74292, 4.74149, 
    4.74005, 4.73861, 4.73718, 4.73574, 4.73452, 4.7334, 4.73228, 4.73117, 
    4.73005, 4.72893, 4.72781, 4.7267, 4.72558, 4.72446, 4.72334, 4.72244, 
    4.7216, 4.72075, 4.71991, 4.71906, 4.71822, 4.71737, 4.71653, 4.71568, 
    4.71484, 4.71399, 4.71315, 4.71239, 4.71177, 4.71116, 4.71055, 4.70993, 
    4.70932, 4.70871, 4.70809, 4.70748, 4.70687, 4.70625, 4.70564, 4.70503, 
    4.70441, 4.7038, 4.70335, 4.70293, 4.70251, 4.70209, 4.70166, 4.70124, 
    4.70082, 4.7004, 4.69998, 4.69956, 4.69913, 4.69871, 4.69829, 4.69787, 
    4.69745, 4.69703, 4.6966, 4.69625, 4.69598, 4.69571, 4.69545, 4.69518, 
    4.69491, 4.69464, 4.69438, 4.69411, 4.69384, 4.69358, 4.69331, 4.69304, 
    4.69278, 4.69251, 4.69224, 4.69197, 4.69171, 4.69144, 4.69117, 4.69091, 
    4.69064, 4.69044, 4.69029, 4.69014, 4.69, 4.68985, 4.6897, 4.68955, 
    4.6894, 4.68925, 4.6891, 4.68895, 4.6888, 4.68866, 4.68851, 4.68836, 
    4.68821, 4.68806, 4.68791, 4.68776, 4.68761, 4.68746, 4.68732, 4.68717, 
    4.68702, 4.68687, 4.68672, 4.68657, 4.68642, 4.68627, 4.68616, 4.68609, 
    4.68603, 4.68596, 4.6859, 4.68583, 4.68577, 4.6857, 4.68563, 4.68557, 
    4.6855, 4.68544, 4.68537, 4.68531, 4.68524, 4.68518, 4.68511, 4.68505, 
    4.68498, 4.68492, 4.68485, 4.68479, 4.68472, 4.68466, 4.68459, 4.68453, 
    4.68446, 4.6844, 4.68433, 4.68427, 4.6842, 4.68414, 4.68407, 4.68401, 
    4.68394, 4.68388, 4.68381, 4.68375, 4.68368, 4.68362, 4.68355, 4.68349, 
    4.68342, 4.68336, 4.68329 ;

 idx_rfr_Fe2O3_doccd_img = 0.04682, 0.04923, 0.05178, 0.05447, 0.0573, 0.0603, 
    0.06346, 0.06681, 0.07035, 0.07408, 0.07805, 0.08224, 0.08668, 0.0914, 
    0.09639, 0.10169, 0.10731, 0.11328, 0.11962, 0.12636, 0.13353, 0.14115, 
    0.14925, 0.15788, 0.16706, 0.17683, 0.18723, 0.1983, 0.21008, 0.22262, 
    0.23595, 0.25011, 0.26516, 0.28112, 0.29803, 0.31592, 0.33481, 0.35472, 
    0.37564, 0.39757, 0.42048, 0.44431, 0.46904, 0.49456, 0.52077, 0.54757, 
    0.57481, 0.60236, 0.63006, 0.65774, 0.68522, 0.71233, 0.73889, 0.76473, 
    0.78968, 0.81358, 0.83627, 0.85762, 0.87751, 0.89583, 0.91248, 0.92741, 
    0.94056, 0.95194, 0.96154, 0.9694, 0.9756, 0.98021, 0.98337, 0.98522, 
    0.98592, 0.98565, 0.98463, 0.98305, 0.98112, 0.97907, 0.97709, 0.97539, 
    0.97414, 0.97348, 0.97355, 0.97439, 0.97604, 0.97845, 0.98148, 0.98497, 
    0.98862, 0.9921, 0.99503, 0.99698, 0.99756, 0.99646, 0.99343, 0.98846, 
    0.98165, 0.97338, 0.96423, 0.95509, 0.94727, 0.94294, 0.94599, 0.96033, 
    0.96066, 0.91959, 0.89362, 0.88579, 0.88707, 0.89418, 0.90609, 0.92243, 
    0.94301, 0.96763, 0.99596, 1.0275, 1.06153, 1.09707, 1.13286, 1.16744, 
    1.19909, 1.22605, 1.24657, 1.25912, 1.26253, 1.2562, 1.24021, 1.21527, 
    1.18272, 1.1443, 1.10205, 1.05801, 1.01412, 0.97213, 0.93352, 0.89959, 
    0.87128, 0.84922, 0.83326, 0.82203, 0.81222, 0.79855, 0.77537, 0.73997, 
    0.69445, 0.64419, 0.59458, 0.54895, 0.50859, 0.4735, 0.44314, 0.41677, 
    0.39374, 0.37344, 0.35541, 0.33926, 0.32469, 0.31146, 0.29937, 0.28827, 
    0.27801, 0.26852, 0.25968, 0.25142, 0.24369, 0.23644, 0.2296, 0.22315, 
    0.21705, 0.21127, 0.20579, 0.20057, 0.1956, 0.19085, 0.18633, 0.182, 
    0.17785, 0.17387, 0.17005, 0.16638, 0.16285, 0.15945, 0.15618, 0.15302, 
    0.14998, 0.14703, 0.14418, 0.14143, 0.13877, 0.13619, 0.13368, 0.13126, 
    0.12891, 0.12662, 0.1244, 0.12225, 0.12015, 0.11811, 0.11612, 0.11419, 
    0.1123, 0.11046, 0.10868, 0.10693, 0.10522, 0.10356, 0.10193, 0.10035, 
    0.0988, 0.09729, 0.09581, 0.09436, 0.09295, 0.09156, 0.09021, 0.08887, 
    0.08757, 0.0863, 0.08505, 0.08383, 0.08263, 0.08146, 0.08031, 0.07918, 
    0.07807, 0.07699, 0.07592, 0.07487, 0.07384, 0.07283, 0.07185, 0.07087, 
    0.06992, 0.06897, 0.06805, 0.06715, 0.06626, 0.06538, 0.06452, 0.06368, 
    0.06284, 0.06202, 0.06122, 0.06043, 0.05964, 0.05888, 0.05813, 0.05738, 
    0.05665, 0.05593, 0.05522, 0.05453, 0.05384, 0.05316, 0.0525, 0.05184, 
    0.0512, 0.05056, 0.04993, 0.04931, 0.04871, 0.0481, 0.04751, 0.04693, 
    0.04636, 0.04579, 0.04524, 0.04469, 0.04415, 0.04362, 0.04309, 0.04257, 
    0.04206, 0.04155, 0.04106, 0.04057, 0.04009, 0.03961, 0.03914, 0.03868, 
    0.03822, 0.03777, 0.03733, 0.03689, 0.03646, 0.03603, 0.03561, 0.0352, 
    0.03479, 0.03439, 0.03399, 0.03359, 0.03321, 0.03283, 0.03245, 0.03208, 
    0.03172, 0.03136, 0.031, 0.03065, 0.0303, 0.02996, 0.02963, 0.0293, 
    0.02897, 0.02865, 0.02833, 0.02802, 0.02771, 0.02741, 0.02711, 0.02681, 
    0.02652, 0.02623, 0.02595, 0.02567, 0.02539, 0.02513, 0.02485, 0.02459, 
    0.02434, 0.02408, 0.02383, 0.02359, 0.02334, 0.02311, 0.02288, 0.02263, 
    0.02241, 0.02219, 0.02197, 0.02175, 0.02154, 0.02133, 0.02112, 0.02093, 
    0.02073, 0.02054, 0.02035, 0.02017, 0.01998, 0.0198, 0.01964, 0.01946, 
    0.0193, 0.01914, 0.01898, 0.01882, 0.01867, 0.01853, 0.01839, 0.01825, 
    0.01812, 0.018, 0.01787, 0.01775, 0.01764, 0.01752, 0.01742, 0.01732, 
    0.01722, 0.01713, 0.01705, 0.01697, 0.01689, 0.01682, 0.01676, 0.01671, 
    0.01665, 0.01661, 0.01657, 0.01654, 0.01651, 0.01649, 0.01649, 0.01648, 
    0.01649, 0.0165, 0.01652, 0.01656, 0.0166, 0.01665, 0.01671, 0.01678, 
    0.01687, 0.01696, 0.01707, 0.01719, 0.01733, 0.01748, 0.01765, 0.01783, 
    0.01803, 0.01825, 0.01849, 0.01876, 0.01903, 0.01934, 0.01968, 0.02005, 
    0.02044, 0.02086, 0.02132, 0.02182, 0.02235, 0.02293, 0.02356, 0.02424, 
    0.02498, 0.02578, 0.02664, 0.02758, 0.0286, 0.02972, 0.03093, 0.03226, 
    0.03371, 0.0353, 0.03706, 0.03899, 0.04114, 0.0435, 0.04617, 0.04914, 
    0.05247, 0.05629, 0.06061, 0.06554, 0.07136, 0.07815, 0.08616, 0.09586, 
    0.10804, 0.12344, 0.14361, 0.1713, 0.21351, 0.2858, 0.41017, 0.58569, 
    0.77339, 0.94991, 1.11444, 1.27086, 1.42264, 1.57267, 1.72345, 1.87715, 
    2.03593, 2.20221, 2.37881, 2.56916, 2.77744, 3.00864, 3.26756, 3.55519, 
    3.84995, 4.0298, 3.8044, 3.13433, 2.43433, 1.9829, 1.83933, 1.95252, 
    2.25645, 2.65018, 3.06164, 3.49079, 3.94823, 4.44823, 5.01553, 5.66556, 
    6.22049, 6.27598, 5.46094, 3.73457, 2.51767, 1.70728, 1.25349, 1.02056, 
    0.85798, 0.75149, 0.69739, 0.67252, 0.6704, 0.70273, 0.78425, 0.91244, 
    1.15604, 1.49635, 1.89202, 2.29379, 2.6838, 3.05941, 3.42943, 3.80023, 
    4.18382, 4.58417, 5.00608, 5.47639, 5.96745, 6.56685, 7.19783, 8.00199, 
    8.88301, 9.97236, 10.90026, 11.56607, 10.72978, 8.06466, 5.77562, 
    3.89923, 2.58499, 1.93947, 1.43985, 1.16981, 0.93594, 0.79989, 0.66961, 
    0.59217, 0.51473, 0.4635, 0.41615, 0.37996, 0.35168, 0.33292, 0.34471, 
    0.35649, 0.32484, 0.28395, 0.24636, 0.2151, 0.18384, 0.16977, 0.16032, 
    0.15124, 0.1442, 0.13715, 0.13074, 0.12516, 0.11957, 0.11467, 0.11016, 
    0.10565, 0.10175, 0.09805, 0.09436, 0.09115, 0.0881, 0.08505, 0.08233, 
    0.0798, 0.07726, 0.0749, 0.07276, 0.07063, 0.06852, 0.06672, 0.06492, 
    0.06312, 0.06148, 0.05995, 0.05842, 0.05689, 0.05558, 0.05426, 0.05295, 
    0.05168, 0.05055, 0.04943, 0.0483, 0.04722, 0.04625, 0.04528, 0.04431, 
    0.04336, 0.04252, 0.04168, 0.04083, 0.03999, 0.03924, 0.03851, 0.03777, 
    0.03704, 0.03634, 0.0357, 0.03507, 0.03444, 0.03381, 0.0332, 0.03265, 
    0.03209, 0.03153, 0.03097, 0.03044, 0.02995, 0.02946, 0.02898, 0.02849, 
    0.02801, 0.02757, 0.02715, 0.02673, 0.0263, 0.02588, 0.02546, 0.02509, 
    0.02472, 0.02435, 0.02398, 0.02362, 0.02325, 0.02291, 0.02259, 0.02226, 
    0.02194, 0.02161, 0.02128, 0.02096, 0.02068, 0.0204, 0.02012, 0.01983, 
    0.01955, 0.01927, 0.01898, 0.01874, 0.01849, 0.01825, 0.018, 0.01776, 
    0.01751, 0.01727, 0.01703, 0.01681, 0.0166, 0.01638, 0.01617, 0.01595, 
    0.01574, 0.01552, 0.01531, 0.0151, 0.01492, 0.01473, 0.01455, 0.01437, 
    0.01418, 0.014, 0.01382, 0.01363, 0.01345, 0.01329, 0.01313, 0.01297, 
    0.01281, 0.01266, 0.0125, 0.01234, 0.01218, 0.01203, 0.01187, 0.01171, 
    0.01157, 0.01144, 0.0113, 0.01117, 0.01104, 0.0109, 0.01077, 0.01063, 
    0.0105, 0.01036, 0.01023, 0.0101, 0.00997, 0.00986, 0.00975, 0.00964, 
    0.00953, 0.00942, 0.0093, 0.00919, 0.00908, 0.00897, 0.00886, 0.00875, 
    0.00864, 0.00853, 0.00842, 0.00832, 0.00823, 0.00813, 0.00804, 0.00795, 
    0.00785, 0.00776, 0.00767, 0.00757, 0.00748, 0.00739, 0.00729, 0.0072, 
    0.0071, 0.00701, 0.00692, 0.00682, 0.00674, 0.00667, 0.0066, 0.00653, 
    0.00646, 0.00639, 0.00633, 0.00626, 0.00619, 0.00612, 0.00605, 0.00598, 
    0.00591, 0.00584, 0.00577, 0.0057, 0.00563, 0.00556, 0.0055, 0.00543, 
    0.00536, 0.00529, 0.00523, 0.00518, 0.00513, 0.00508, 0.00503, 0.00498, 
    0.00493, 0.00488, 0.00482, 0.00477, 0.00472, 0.00467, 0.00462, 0.00457, 
    0.00452, 0.00447, 0.00442, 0.00437, 0.00432, 0.00427, 0.00422, 0.00417, 
    0.00412, 0.00407, 0.00401, 0.00396, 0.00391, 0.00386, 0.00381, 0.00377, 
    0.00373, 0.00369, 0.00366, 0.00362, 0.00359, 0.00355, 0.00351, 0.00348, 
    0.00344, 0.00341, 0.00337, 0.00333, 0.0033, 0.00326, 0.00323, 0.00319, 
    0.00315, 0.00312, 0.00308, 0.00305, 0.00301, 0.00297, 0.00294, 0.0029, 
    0.00287, 0.00283, 0.00279, 0.00276, 0.00272, 0.00268, 0.00265, 0.00261, 
    0.00258, 0.00254, 0.0025, 0.00247, 0.00243, 0.0024, 0.00236, 0.00232, 
    0.00229, 0.00225, 0.00222, 0.00218 ;
}

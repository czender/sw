// $Id$
// ncgen -b -o ${DATA}/aca/idx_rfr_shettle_Fe2O3_SiO2.nc ${HOME}/idx_rfr/idx_rfr_shettle_Fe2O3_SiO2.cdl
// Define "_avg" indices of refraction as average of O-ray and E-ray indices
// ncap -O -s 'idx_rfr_Fe2O3_avg_hitran96_rl=0.5*(idx_rfr_Fe2O3_oray_hitran96_rl+idx_rfr_Fe2O3_eray_hitran96_rl)' -s 'idx_rfr_Fe2O3_avg_hitran96_img=0.5*(idx_rfr_Fe2O3_oray_hitran96_img+idx_rfr_Fe2O3_eray_hitran96_img)' -s 'idx_rfr_SiO2_avg_hitran96_rl=0.5*(idx_rfr_SiO2_oray_hitran96_rl+idx_rfr_SiO2_eray_hitran96_rl)' -s 'idx_rfr_SiO2_avg_hitran96_img=0.5*(idx_rfr_SiO2_oray_hitran96_img+idx_rfr_SiO2_eray_hitran96_img)' ${DATA}/aca/idx_rfr_shettle_Fe2O3_SiO2.nc ${DATA}/aca/idx_rfr_shettle_Fe2O3_SiO2.nc

netcdf idx_rfr_shettle_Fe2O3_SiO2 {
dimensions:
	bnd=68;
variables:

	:RCS_Header = "$Id$";
	:history = "";
	:source="HITRAN96 CDROM file /cdrom/aerosols/shettle.dat,
Table A5
Standardized by Charlie Zender 20041226
		   TABLE A5
  ---------------------------------------------------                                                                                
 Quartz            A-15, A-16, A-17,  Anisotropic material. 
                   A-18, A-19         Values are given for  
                                      the O and E rays      
                                                            
 Hematite          A-19, A-20, A-21,  Anisotropic material. 
 (Iron Oxide)      A-22, A-23         Values are given for  
                                      the O and E rays      
 ----------------------------------------------------                                    
A-15. Gray, D. C. (1963), American Institute of Physics Handbook,
McGraw-Hill, New York, NY, 1963, 2nd Edition.

A-16. Drummond, D. G. (1936) Absorption coefficients of crystal
quartz in the infrared, Proc. Roy. Soc. (London)-Series A,
153:328-338.

A-17. Spitzer, W. G. and Kleinman, D. A. (1961) Infrared lattice
bands of quartz, Phys. Rev., 121:1324-1335.

A-18. Philipp, H. R. (1985) Silicon dioxide (SiO2), type-
(crystalline), in Handbook of Optical Constants of Solids, Edited
by E. D. Palik, Academic Press, Inc., Orlando, FL, 719-747.

A-19. Longtin, D. R., Shettle, E. P., Hummel, J. R. and Pryce, J.
D., (1988) A Wind Dependent Desert Aerosol Model: Radiative
Properties, AFGL-TR-88-0112, Air Force Geophysics Laboratory,
Hanscom AFB, MA, April 1988.

A-20. Galuza, A. I., Eremenko, V. V. and Kirichenko, A. P. (1979)
Analysis of hematite reflection spectrum by the Kramers-Kronig
method, Sov. Phys. Solid State, 21:654-656.

A-21. Kerker, M., Scheiner, P., Cooke, D. D. and Kratohvil, J.P.
(1979) Absorption index and color of colloidal hematite, J.
Colloid. Interface Sci., 71:176-187.

A-22. Steyer, T. R. (1974) Infrared optical properties of some
solids of possible interest in astronomy and atmospheric physics,
Graduate Thesis, Department of Physics, University of Arizona.

A-23. Onari, S., Arai, T. and Kudo, K. (1977) Infrared lattice
vibrations and dielectric dispersion in - Fe2O3, Phys. Rev. B,
16:1717-1721.";

	float bnd(bnd);
	bnd:long_name = "Band center wavelength";
	bnd:units = "micron";
	bnd:C_format = "%.5g";

	float idx_rfr_Fe2O3_oray_hitran96_rl(bnd);
	idx_rfr_Fe2O3_oray_hitran96_rl:long_name = "Hematite real index of refraction O-ray";
	idx_rfr_Fe2O3_oray_hitran96_rl:units = "";
	idx_rfr_Fe2O3_oray_hitran96_rl:composition = "Fe2O3";
	idx_rfr_Fe2O3_oray_hitran96_rl:C_format = "%.4g";

	float idx_rfr_Fe2O3_oray_hitran96_img(bnd);
	idx_rfr_Fe2O3_oray_hitran96_img:long_name = "Hematite imaginary index of refraction O-ray";
	idx_rfr_Fe2O3_oray_hitran96_img:units = "";
	idx_rfr_Fe2O3_oray_hitran96_img:composition = "Fe2O3";
	idx_rfr_Fe2O3_oray_hitran96_img:C_format = "%.3g";

	float idx_rfr_Fe2O3_eray_hitran96_rl(bnd);
	idx_rfr_Fe2O3_eray_hitran96_rl:long_name = "Hematite real index of refraction E-ray";
	idx_rfr_Fe2O3_eray_hitran96_rl:units = "";
	idx_rfr_Fe2O3_eray_hitran96_rl:composition = "Fe2O3";
	idx_rfr_Fe2O3_eray_hitran96_rl:C_format = "%.4g";

	float idx_rfr_Fe2O3_eray_hitran96_img(bnd);
	idx_rfr_Fe2O3_eray_hitran96_img:long_name = "Hematite imaginary index of refraction E-ray";
	idx_rfr_Fe2O3_eray_hitran96_img:units = "";
	idx_rfr_Fe2O3_eray_hitran96_img:composition = "Fe2O3";
	idx_rfr_Fe2O3_eray_hitran96_img:C_format = "%.3g";

	float idx_rfr_SiO2_oray_hitran96_rl(bnd);
	idx_rfr_SiO2_oray_hitran96_rl:long_name = "Quartz real index of refraction O-ray";
	idx_rfr_SiO2_oray_hitran96_rl:units = "";
	idx_rfr_SiO2_oray_hitran96_rl:composition = "SiO2";
	idx_rfr_SiO2_oray_hitran96_rl:C_format = "%.4g";

	float idx_rfr_SiO2_oray_hitran96_img(bnd);
	idx_rfr_SiO2_oray_hitran96_img:long_name = "Quartz imaginary index of refraction O-ray";
	idx_rfr_SiO2_oray_hitran96_img:units = "";
	idx_rfr_SiO2_oray_hitran96_img:composition = "SiO2";
	idx_rfr_SiO2_oray_hitran96_img:C_format = "%.3g";

	float idx_rfr_SiO2_eray_hitran96_rl(bnd);
	idx_rfr_SiO2_eray_hitran96_rl:long_name = "Quartz real index of refraction E-ray";
	idx_rfr_SiO2_eray_hitran96_rl:units = "";
	idx_rfr_SiO2_eray_hitran96_rl:composition = "SiO2";
	idx_rfr_SiO2_eray_hitran96_rl:C_format = "%.4g";

	float idx_rfr_SiO2_eray_hitran96_img(bnd);
	idx_rfr_SiO2_eray_hitran96_img:long_name = "Quartz imaginary index of refraction E-ray";
	idx_rfr_SiO2_eray_hitran96_img:units = "";
	idx_rfr_SiO2_eray_hitran96_img:composition = "SiO2";
	idx_rfr_SiO2_eray_hitran96_img:C_format = "%.3g";

data:	
 bnd =    0.200,   0.250,   0.300,   0.337,   0.400,
   0.488,   0.515,   0.550,   0.633,   0.694,
   0.860,   1.060,   1.300,   1.536,   1.800,
   2.000,   2.250,   2.500,   2.700,   3.000,
   3.200,   3.392,   3.500,   3.750,   4.000,
   4.500,   5.000,   5.500,   6.000,   6.200,
   6.500,   7.200,   7.900,   8.200,   8.500,
   8.700,   9.000,   9.200,   9.500,   9.800,
  10.000,  10.591,  11.000,  11.500,  12.500,
  13.000,  14.000,  14.800,  15.000,  16.400,
  17.200,  18.000,  18.500,  20.000,  21.300,
  22.500,  25.000,  27.900,  30.000,  35.000,
  40.000,  50.000,  60.000,  80.000, 100.000,
 150.000, 200.000, 300.000;
 
 idx_rfr_SiO2_oray_hitran96_rl = 1.649,1.606,1.584,1.568,1.559,
1.550,1.548,1.546,1.542,1.541,
1.537,1.534,1.531,1.538,1.524,
1.520,1.516,1.511,1.506,1.499,
1.493,1.487,1.483,1.473,1.462,
1.442,1.417,1.371,1.325,1.293,
1.246,1.065,0.585,0.141,0.114,
0.131,0.176,0.633,4.497,3.014,
2.663,2.188,2.013,1.833,1.587,
2.174,1.768,1.831,1.785,1.580,
1.456,1.289,1.142,0.106,0.194,
5.709,0.679,2.729,2.500,2.305,
2.228,2.214,2.175,2.148,2.132,
2.120,2.111,2.109;

 idx_rfr_SiO2_oray_hitran96_img = 1.0e-8 ,1.0e-8 ,1.0e-8 ,1.0e-8 ,1.0e-8 ,
1.0e-8 ,1.0e-8 ,1.0e-8 ,1.0e-8 ,1.0e-8 ,
1.0e-8 ,1.0e-8 ,1.0e-8 ,1.0e-8 ,1.0e-8 ,
1.0e-8 ,1.0e-8 ,4.99e-7,7.20e-7,2.67e-5,
6.77e-6,6.40e-6,8.31e-6,5.95e-5,7.12e-5,
5.06e-4,0.00562,0.00551,0.00674,0.00782,
0.00580,0.0124 ,0.0849 ,0.538  ,1.26   ,
1.41   ,2.61   ,4.55   ,0.392  ,0.0869 ,
0.0517 ,0.0222 ,0.0173 ,0.0188 ,2.27   ,
0.0519 ,0.0348 ,0.0229 ,0.0154 ,0.00975,
0.0120 ,0.0177 ,0.0252 ,0.766  ,2.57   ,
0.941  ,1.85   ,0.0216 ,0.0108 ,0.00498,
0.00329,0.00286,0.00224,0.00369,9.55e-4,
8.72e-4,7.96e-4,7.96e-4;

 idx_rfr_SiO2_eray_hitran96_rl = 1.649,1.606,1.584,1.568,1.559,
1.550,1.548,1.546,1.542,1.541,
1.537,1.534,1.531,1.528,1.524,
1.520,1.516,1.511,1.506,1.499,
1.493,1.487,1.483,1.473,1.462,
1.442,1.417,1.371,1.325,1.293,
1.246,1.063,0.564,0.123,0.085,
0.096,0.231,1.689,3.899,2.860,
2.571,2.156,1.999,1.849,1.260,
2.625,1.821,1.670,1.636,1.361,
1.093,0.425,0.197,1.270,3.041,
2.366,1.451,4.905,2.959,2.464,
2.337,2.262,2.223,2.190,2.176,
2.163,2.159,2.156;

 idx_rfr_SiO2_eray_hitran96_img = 1.0e-8 ,1.0e-8 ,1.0e-8 ,1.0e-8 ,1.0e-8 ,
1.0e-8 ,1.0e-8 ,1.0e-8 ,1.0e-8 ,1.0e-8 ,
1.0e-8 ,1.0e-8 ,1.0e-8 ,1.0e-8 ,1.0e-8 ,
1.0e-8 ,1.0e-8 ,7.48e-7,1.14e-6,8.47e-6,
4.03e-6,5.70e-6,8.31e-6,3.68e-5,7.12e-5,
3.58e-4,0.00446,0.00520,0.00480,0.00782,
0.00730,0.0146 ,0.0861 ,0.586  ,1.22   ,
1.72   ,3.05   ,6.41   ,0.229  ,0.0691 ,
0.0440 ,0.0205 ,0.0159 ,0.0153 ,0.130  ,
0.318  ,0.0165 ,0.0121 ,0.0121 ,0.0192 ,
0.0377 ,0.212  ,0.973  ,4.98   ,0.102  ,
0.0438 ,0.0999 ,0.860  ,0.0593 ,0.0125 ,
0.00675,0.00171,0.00108,6.35e-4,4.77e-4,
2.40e-4,1.59e-4,6.20e-5;

 idx_rfr_Fe2O3_oray_hitran96_rl = 1.560,2.070,2.320,2.430,2.674,
3.074,3.104,3.102,3.007,2.920,
2.730,2.690,2.660,2.640,2.620,
2.610,2.610,2.610,2.610,2.610,
2.610,2.610,2.610,2.610,2.670,
2.660,2.650,2.640,2.620,2.610,
2.590,2.540,2.490,2.450,2.420,
2.400,2.370,2.340,2.300,2.260,
2.240,2.140,2.069,1.970,1.760,
1.645,1.225,0.742,0.554,0.194,
0.265,0.520,1.097,2.042,0.941,
3.306,3.714,0.591,0.430,15.362,
7.621,6.349,5.671,5.266,5.122,
4.998,4.958,4.931;

 idx_rfr_Fe2O3_oray_hitran96_img = 1.28   ,1.33   ,1.18   ,1.09   ,0.523  ,
0.210  ,0.158  ,0.0925 ,0.00974,0.00100,
0.00400,3.0e-5 ,1.8e-5 ,1.3e-5 ,1.1e-5 ,
1.0e-5 ,1.0e-5 ,1.0e-5 ,1.0e-5 ,1.0e-5 ,
1.1e-5 ,1.1e-5 ,1.2e-5 ,1.2e-5 ,6.7e-5 ,
6.0e-5 ,5.3e-5 ,6.2e-4 ,0.0012 ,0.0015 ,
0.0017 ,0.0018 ,0.0018 ,0.0031 ,0.0044 ,
0.0057 ,0.0070 ,0.0076 ,0.0085 ,0.0094 ,
0.0100 ,0.0145 ,0.0174 ,0.0216 ,0.0367 ,
0.0477 ,0.0675 ,0.204  ,0.295  ,1.56   ,
2.25   ,3.13   ,3.89   ,1.63   ,3.61   ,
6.22   ,0.684  ,2.06   ,4.31   ,13.9   ,
0.387  ,0.107  ,0.0533 ,0.0290 ,0.0205 ,
0.0122 ,0.00886,0.00576;

 idx_rfr_Fe2O3_eray_hitran96_rl = 1.560,2.070,2.320,2.430,2.674,
3.074,3.104,3.102,3.007,2.920,
2.730,2.690,2.660,2.640,2.620,
2.610,2.610,2.610,2.610,2.610,
2.610,2.610,2.610,2.610,2.470,
2.460,2.440,2.420,2.400,2.390,
2.380,2.340,2.300,2.270,2.250,
2.230,2.210,2.190,2.160,2.130,
2.110,2.031,1.972,1.894,1.720,
1.618,1.286,0.823,0.668,0.343,
0.519,1.093,2.212,4.351,3.048,
2.209,0.520,0.492,0.889,10.861,
6.869,5.479,5.080,4.792,4.683,
4.587,4.555,4.534; 

 idx_rfr_Fe2O3_eray_hitran96_img = 1.28   ,1.33   ,1.18   ,1.09   ,0.523  ,
0.210  ,0.158  ,0.0925 ,0.00974,0.00100,
0.00400,3.0e-5 ,1.8e-5 ,1.3e-5 ,1.1e-5 ,
1.0e-5 ,1.0e-5 ,1.0e-5 ,1.0e-5 ,1.0e-5 ,
1.1e-5 ,1.1e-5 ,1.2e-5 ,1.2e-5 ,1.3e-5 ,
1.9e-5 ,2.5e-5 ,3.0e-5 ,3.5e-5 ,3.4e-5 ,
3.2e-5 ,6.0e-5 ,8.0e-5 ,3.0e-4 ,5.0e-4 ,
8.0e-4 ,0.0010 ,0.0026 ,0.0050 ,0.0074 ,
0.0090 ,0.0126 ,0.0151 ,0.0207 ,0.0364 ,
0.0472 ,0.105  ,0.243  ,0.331  ,1.79   ,
2.64   ,3.78   ,4.65   ,1.14   ,0.487  ,
0.417  ,1.69   ,3.91   ,5.95   ,2.58   ,
0.388  ,0.121  ,0.0713 ,0.0404 ,0.0289 ,
0.0173 ,0.0125 ,0.00816;

}

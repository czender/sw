// $Id$
// ncgen -b -o ${DATA}/aca/idx_rfr_Fe2O3.nc ${HOME}/idx_rfr/idx_rfr_Fe2O3.cdl
// Define "_avg" indices of refraction as average of O-ray and E-ray indices
// ncap -O -s 'idx_rfr_Fe2O3_avg_roush_rl=0.5*(idx_rfr_Fe2O3_oray_roush_rl+idx_rfr_Fe2O3_eray_roush_rl)' -s 'idx_rfr_Fe2O3_avg_roush_img=0.5*(idx_rfr_Fe2O3_oray_roush_img+idx_rfr_Fe2O3_eray_roush_img)' ${DATA}/aca/idx_rfr_Fe2O3.nc ${DATA}/aca/idx_rfr_Fe2O3.nc
// rsync ${DATA}/aca/idx_rfr_Fe2O3.nc esmf.ess.uci.edu:/data/zender/aca

netcdf idx_rfr_Fe2O3 {
dimensions:
	bnd = 613 ;

variables:

// global attributes:
	:RCS_Header = "$Id$" ;
	:history = "" ;
	:description = "Hematite refractive indices" ;
	:source="
Ted Roush (NASA Ames) <troush at mail dot arc dot nasa dot gov>
Charlie Zender (UCI) <zender at uci dot edu> standardized 20060630.

Changes:
Changed coordinate from wavenumber to wavelength.
Extended data from 0.21 um to 0.20 um by copying 0.21 um data.
Took absolute value of four negative imaginary refractive indices near 50 um.

Begin Procedure to create netCDF from text file:
fl_txt=idx_rfr_Fe2O3
cat > /tmp/${fl_txt}.header << EOF
bnd_wvn_Fe2O3_oray_roush:f bnd:f idx_rfr_Fe2O3_oray_roush_rl:f idx_rfr_Fe2O3_oray_roush_img:f idx_rfr_Fe2O3_oray_roush_rl_ee:f idx_rfr_Fe2O3_oray_roush_img_ee:f idx_rfr_Fe2O3_oray_roush_nr:f
EOF
tbl2cdf -h /tmp/${fl_txt}.header ~/hematite.txt ~/idx_rfr/${fl_txt}.nc
ncrename -O -d u,bnd ${fl_txt}.nc
ncks ~/idx_rfr/${fl_txt}.nc | m
ncdump ~/idx_rfr/${fl_txt}.nc > ~/${fl_txt}.cdl
End Procedure to create netCDF from text file:

Begin Original e-mail header accompanying data from T. Roush:
From:	IO::memilham@CRDEC-VAX4.ARPA 14-JUN-1988 12:56
To:	HAL::DALTON
Subj:	Optical Constants: Hematite E-Ray

Received: from CRDEC-VAX4.ARPA by ames-io.ARPA with INTERNET ;
          Tue, 14 Jun 88 12:44:14 PDT
Date:     Tue, 14 Jun 88 14:23:02 EDT
From:     Merrill E. Milham <memilham@CRDEC-VAX4.ARPA>
To:       dalton%hal@AMES-IO.ARPA
Subject:  Optical Constants: Hematite E-Ray
Message-ID:  <8806141423.aa16177@CRDEC-VAX4.CRDEC-VAX4.ARPA>
 
HEMITE E-RAY M.R.QUERRY
        wn     wl        n       k      Dn       Dk      R
       (cm-1) (um)

From:	IO::memilham@CRDEC-VAX4.ARPA 14-JUN-1988 12:53
To:	HAL::DALTON
Subj:	Optical Constants: Hematite O-Ray

Received: from CRDEC-VAX4.ARPA by ames-io.ARPA with INTERNET ;
          Tue, 14 Jun 88 12:43:20 PDT
Date:     Tue, 14 Jun 88 14:21:25 EDT
From:     Merrill E. Milham <memilham@CRDEC-VAX4.ARPA>
To:       dalton%hal@AMES-IO.ARPA
Subject:  Optical Constants: Hematite O-Ray
Message-ID:  <8806141421.aa16102@CRDEC-VAX4.CRDEC-VAX4.ARPA>
 
HEMATITE O-RAY  M.R.QUERRY
        wn      wl       n       k       Dn      Dk      R
       (cm-1)  (um)
End Original e-mail header accompanying data from T. Roush
	";

	float bnd(bnd) ;
		bnd:units = "microns" ;
		bnd:longname = "Band center wavelength" ;
		bnd:C_format = "%.5g" ;

	float bnd_wvn_Fe2O3_eray_roush(bnd) ;
		bnd_wvn_Fe2O3_eray_roush:units = "cm-1" ;
		bnd_wvn_Fe2O3_eray_roush:longname = "Band center wavenumber" ;
		bnd_wvn_Fe2O3_eray_roush:C_format = "%.5g" ;

	float idx_rfr_Fe2O3_eray_roush_rl(bnd) ;
		idx_rfr_Fe2O3_eray_roush_rl:units = "" ;
		idx_rfr_Fe2O3_eray_roush_rl:longname = "Hematite refractive index, real part, E-ray" ;
		idx_rfr_Fe2O3_eray_roush_rl:C_format = "%.4g" ;

	float idx_rfr_Fe2O3_eray_roush_img(bnd) ;
		idx_rfr_Fe2O3_eray_roush_img:units = "" ;
		idx_rfr_Fe2O3_eray_roush_img:longname = "Hematite refractive index, imaginary part, E-ray" ;
		idx_rfr_Fe2O3_eray_roush_img:C_format = "%.3g" ;

	float idx_rfr_Fe2O3_eray_roush_rl_ee(bnd) ;
		idx_rfr_Fe2O3_eray_roush_rl_ee:units = "" ;
		idx_rfr_Fe2O3_eray_roush_rl_ee:longname = "Hematite refractive index estimated error, real part, E-ray" ;
		idx_rfr_Fe2O3_eray_roush_rl_ee:C_format = "%.4g" ;

	float idx_rfr_Fe2O3_eray_roush_img_ee(bnd) ;
		idx_rfr_Fe2O3_eray_roush_img_ee:units = "" ;
		idx_rfr_Fe2O3_eray_roush_img_ee:longname = "Hematite refractive index estimated error, imaginary part, E-ray" ;
		idx_rfr_Fe2O3_eray_roush_img_ee:C_format = "%.3g" ;

	float idx_rfr_Fe2O3_eray_roush_nr(bnd) ;
		idx_rfr_Fe2O3_eray_roush_nr:units = "" ;
		idx_rfr_Fe2O3_eray_roush_nr:longname = "Hematite measured normal reflectance, E-ray" ;
		idx_rfr_Fe2O3_eray_roush_nr:C_format = "%.3g" ;

	float bnd_wvn_Fe2O3_oray_roush(bnd) ;
		bnd_wvn_Fe2O3_oray_roush:units = "cm-1" ;
		bnd_wvn_Fe2O3_oray_roush:longname = "Band center wavenumber" ;
		bnd_wvn_Fe2O3_oray_roush:C_format = "%.5g" ;

	float idx_rfr_Fe2O3_oray_roush_rl(bnd) ;
		idx_rfr_Fe2O3_oray_roush_rl:units = "" ;
		idx_rfr_Fe2O3_oray_roush_rl:longname = "Hematite refractive index, real part, O-ray" ;
		idx_rfr_Fe2O3_oray_roush_rl:C_format = "%.4g" ;

	float idx_rfr_Fe2O3_oray_roush_img(bnd) ;
		idx_rfr_Fe2O3_oray_roush_img:units = "" ;
		idx_rfr_Fe2O3_oray_roush_img:longname = "Hematite refractive index, imaginary part, O-ray" ;
		idx_rfr_Fe2O3_oray_roush_img:C_format = "%.3g" ;

	float idx_rfr_Fe2O3_oray_roush_rl_ee(bnd) ;
		idx_rfr_Fe2O3_oray_roush_rl_ee:units = "" ;
		idx_rfr_Fe2O3_oray_roush_rl_ee:longname = "Hematite refractive index estimated error, real part, O-ray" ;
		idx_rfr_Fe2O3_oray_roush_rl_ee:C_format = "%.4g" ;

	float idx_rfr_Fe2O3_oray_roush_img_ee(bnd) ;
		idx_rfr_Fe2O3_oray_roush_img_ee:units = "" ;
		idx_rfr_Fe2O3_oray_roush_img_ee:longname = "Hematite refractive index estimated error, imaginary part, O-ray" ;
		idx_rfr_Fe2O3_oray_roush_img_ee:C_format = "%.3g" ;

	float idx_rfr_Fe2O3_oray_roush_nr(bnd) ;
		idx_rfr_Fe2O3_oray_roush_nr:units = "" ;
		idx_rfr_Fe2O3_oray_roush_nr:longname = "Hematite measured normal reflectance, O-ray" ;
		idx_rfr_Fe2O3_oray_roush_nr:C_format = "%.3g" ;

data:

 bnd_wvn_Fe2O3_eray_roush = 180, 190, 200, 210, 220, 230, 240, 250, 260, 270, 280, 290, 300, 
    310, 320, 330, 340, 350, 360, 370, 380, 390, 400, 410, 420, 430, 440, 
    450, 460, 470, 480, 490, 500, 510, 520, 530, 540, 550, 560, 570, 580, 
    590, 600, 610, 620, 630, 640, 650, 660, 670, 680, 690, 700, 710, 720, 
    730, 740, 750, 760, 770, 780, 790, 800, 810, 820, 830, 840, 850, 860, 
    870, 880, 890, 900, 910, 920, 930, 940, 950, 960, 970, 980, 990, 1000, 
    1010, 1020, 1030, 1040, 1050, 1060, 1070, 1080, 1090, 1100, 1110, 1120, 
    1130, 1140, 1150, 1160, 1170, 1180, 1190, 1200, 1210, 1220, 1230, 1240, 
    1250, 1260, 1270, 1280, 1290, 1300, 1310, 1320, 1330, 1340, 1350, 1360, 
    1370, 1380, 1390, 1400, 1410, 1420, 1430, 1440, 1450, 1460, 1470, 1480, 
    1490, 1500, 1510, 1520, 1530, 1540, 1550, 1560, 1570, 1580, 1590, 1600, 
    1610, 1620, 1630, 1640, 1650, 1660, 1670, 1680, 1690, 1700, 1710, 1720, 
    1730, 1740, 1750, 1760, 1770, 1780, 1790, 1800, 1810, 1820, 1830, 1840, 
    1850, 1860, 1870, 1880, 1890, 1900, 1910, 1920, 1930, 1940, 1950, 1960, 
    1970, 1980, 1990, 2000, 2010, 2020, 2030, 2040, 2050, 2060, 2070, 2080, 
    2090, 2100, 2110, 2120, 2130, 2140, 2150, 2160, 2170, 2180, 2190, 2200, 
    2210, 2220, 2230, 2240, 2250, 2260, 2270, 2280, 2290, 2300, 2310, 2320, 
    2330, 2340, 2350, 2360, 2370, 2380, 2390, 2400, 2410, 2420, 2430, 2440, 
    2450, 2460, 2470, 2480, 2490, 2500, 2510, 2520, 2530, 2540, 2550, 2560, 
    2570, 2580, 2590, 2600, 2610, 2620, 2630, 2640, 2650, 2660, 2670, 2680, 
    2690, 2700, 2710, 2720, 2730, 2740, 2750, 2760, 2770, 2780, 2790, 2800, 
    2810, 2820, 2830, 2840, 2850, 2860, 2870, 2880, 2890, 2900, 2910, 2920, 
    2930, 2940, 2950, 2960, 2970, 2980, 2990, 3000, 3010, 3020, 3030, 3040, 
    3050, 3060, 3070, 3080, 3090, 3100, 3110, 3120, 3130, 3140, 3150, 3160, 
    3170, 3180, 3190, 3200, 3210, 3220, 3230, 3240, 3250, 3260, 3270, 3280, 
    3290, 3300, 3310, 3320, 3330, 3340, 3350, 3360, 3370, 3380, 3390, 3400, 
    3410, 3420, 3430, 3440, 3450, 3460, 3470, 3480, 3490, 3500, 3510, 3520, 
    3530, 3540, 3550, 3560, 3570, 3580, 3590, 3600, 3610, 3620, 3630, 3640, 
    3650, 3660, 3670, 3680, 3690, 3700, 3710, 3720, 3730, 3740, 3750, 3760, 
    3770, 3780, 3790, 3800, 3810, 3820, 3830, 3840, 3850, 3860, 3870, 3880, 
    3890, 3900, 3910, 3920, 3930, 3940, 3950, 3960, 3970, 3980, 3990, 4000, 
    4016.06, 4032.26, 4048.58, 4065.04, 4081.63, 4098.36, 4115.23, 4132.23, 
    4149.38, 4166.67, 4184.1, 4201.68, 4219.41, 4237.29, 4255.32, 4273.5, 
    4291.85, 4310.34, 4329, 4347.83, 4366.81, 4385.96, 4405.29, 4424.78, 
    4444.44, 4464.29, 4484.3, 4504.5, 4524.89, 4545.45, 4566.21, 4587.16, 
    4608.29, 4629.63, 4651.16, 4672.9, 4694.84, 4716.98, 4739.34, 4761.9, 
    4784.69, 4807.69, 4830.92, 4854.37, 4878.05, 4901.96, 4926.11, 4950.5, 
    4975.12, 5000, 5025.13, 5050.51, 5076.14, 5102.04, 5128.21, 5154.64, 
    5181.35, 5208.33, 5235.6, 5263.16, 5291.01, 5319.15, 5347.59, 5376.34, 
    5405.41, 5434.78, 5464.48, 5494.51, 5524.86, 5555.56, 5586.59, 5617.98, 
    5649.72, 5681.82, 5714.29, 5747.13, 5780.35, 5813.95, 5847.95, 5882.35, 
    5917.16, 5952.38, 5988.02, 6024.1, 6060.61, 6097.56, 6134.97, 6172.84, 
    6211.18, 6250, 6289.31, 6329.11, 6369.43, 6410.26, 6451.61, 6493.51, 
    6535.95, 6578.95, 6622.52, 6666.67, 6711.41, 6756.76, 6802.72, 6849.32, 
    6896.55, 6944.44, 6993.01, 7042.25, 7092.2, 7142.86, 7194.24, 7246.38, 
    7299.27, 7352.94, 7407.41, 7462.69, 7518.8, 7575.76, 7633.59, 7692.31, 
    7751.94, 7812.5, 7874.02, 7936.51, 8000, 8064.52, 8130.08, 8196.72, 
    8264.46, 8333.33, 8403.36, 8474.58, 8547.01, 8620.69, 8695.65, 8771.93, 
    8849.56, 8928.57, 9009.01, 9090.91, 9174.31, 9259.26, 9345.79, 9433.96, 
    9523.81, 9615.38, 9708.74, 9803.92, 9900.99, 10000, 10101.01, 10204.08, 
    10309.28, 10416.67, 10526.32, 10638.3, 10752.69, 10869.57, 10989.01, 
    11111.11, 11235.96, 11363.64, 11494.25, 11627.91, 11764.71, 11904.76, 
    12048.19, 12195.12, 12345.68, 12500, 12658.23, 12820.51, 12987.01, 
    13157.89, 13333.33, 13513.51, 13698.63, 13888.89, 14084.51, 14285.71, 
    14492.75, 14705.88, 14925.37, 15151.52, 15384.62, 15625, 15873.02, 
    16129.03, 16393.44, 16666.67, 16949.15, 17241.38, 17543.86, 17857.14, 
    18181.82, 18518.52, 18867.92, 19230.77, 19607.84, 20000, 20408.16, 
    20833.33, 21276.6, 21739.13, 22222.22, 22727.27, 23255.81, 23809.52, 
    24390.24, 25000, 25641.03, 26315.79, 27027.03, 27777.78, 28571.43, 
    29411.76, 30303.03, 31250, 32258.06, 33333.33, 34482.76, 35714.29, 
    37037.04, 38461.54, 40000, 41666.67, 43478.26, 45454.55, 47619.05,
// Copy data from 0.21 um to 0.20 um
	50000.0 ;

 bnd = 55.5556, 52.6316, 50, 47.619, 45.4545, 43.4783, 41.6667, 40, 38.4615, 
    37.037, 35.7143, 34.4828, 33.3333, 32.2581, 31.25, 30.303, 29.4118, 
    28.5714, 27.7778, 27.027, 26.3158, 25.641, 25, 24.3902, 23.8095, 23.2558, 
    22.7273, 22.2222, 21.7391, 21.2766, 20.8333, 20.4082, 20, 19.6078, 
    19.2308, 18.8679, 18.5185, 18.1818, 17.8571, 17.5439, 17.2414, 16.9492, 
    16.6667, 16.3934, 16.129, 15.873, 15.625, 15.3846, 15.1515, 14.9254, 
    14.7059, 14.4928, 14.2857, 14.0845, 13.8889, 13.6986, 13.5135, 13.3333, 
    13.1579, 12.987, 12.8205, 12.6582, 12.5, 12.3457, 12.1951, 12.0482, 
    11.9048, 11.7647, 11.6279, 11.4943, 11.3636, 11.236, 11.1111, 10.989, 
    10.8696, 10.7527, 10.6383, 10.5263, 10.4167, 10.3093, 10.2041, 10.101, 
    10, 9.901, 9.8039, 9.7087, 9.6154, 9.5238, 9.434, 9.3458, 9.2593, 9.1743, 
    9.0909, 9.009, 8.9286, 8.8496, 8.7719, 8.6957, 8.6207, 8.547, 8.4746, 
    8.4034, 8.3333, 8.2645, 8.1967, 8.1301, 8.0645, 8, 7.9365, 7.874, 7.8125, 
    7.7519, 7.6923, 7.6336, 7.5758, 7.5188, 7.4627, 7.4074, 7.3529, 7.2993, 
    7.2464, 7.1942, 7.1429, 7.0922, 7.0423, 6.993, 6.9444, 6.8966, 6.8493, 
    6.8027, 6.7568, 6.7114, 6.6667, 6.6225, 6.5789, 6.5359, 6.4935, 6.4516, 
    6.4103, 6.3694, 6.3291, 6.2893, 6.25, 6.2112, 6.1728, 6.135, 6.0976, 
    6.0606, 6.0241, 5.988, 5.9524, 5.9172, 5.8824, 5.848, 5.814, 5.7803, 
    5.7471, 5.7143, 5.6818, 5.6497, 5.618, 5.5866, 5.5556, 5.5249, 5.4945, 
    5.4645, 5.4348, 5.4054, 5.3763, 5.3476, 5.3191, 5.291, 5.2632, 5.2356, 
    5.2083, 5.1813, 5.1546, 5.1282, 5.102, 5.0761, 5.0505, 5.0251, 5, 4.9751, 
    4.9505, 4.9261, 4.902, 4.878, 4.8544, 4.8309, 4.8077, 4.7847, 4.7619, 
    4.7393, 4.717, 4.6948, 4.6729, 4.6512, 4.6296, 4.6083, 4.5872, 4.5662, 
    4.5455, 4.5249, 4.5045, 4.4843, 4.4643, 4.4444, 4.4248, 4.4053, 4.386, 
    4.3668, 4.3478, 4.329, 4.3103, 4.2918, 4.2735, 4.2553, 4.2373, 4.2194, 
    4.2017, 4.1841, 4.1667, 4.1494, 4.1322, 4.1152, 4.0984, 4.0816, 4.065, 
    4.0486, 4.0323, 4.0161, 4, 3.9841, 3.9683, 3.9526, 3.937, 3.9216, 3.9063, 
    3.8911, 3.876, 3.861, 3.8462, 3.8314, 3.8168, 3.8023, 3.7879, 3.7736, 
    3.7594, 3.7453, 3.7313, 3.7175, 3.7037, 3.69, 3.6765, 3.663, 3.6496, 
    3.6364, 3.6232, 3.6101, 3.5971, 3.5842, 3.5714, 3.5587, 3.5461, 3.5336, 
    3.5211, 3.5088, 3.4965, 3.4843, 3.4722, 3.4602, 3.4483, 3.4364, 3.4247, 
    3.413, 3.4014, 3.3898, 3.3784, 3.367, 3.3557, 3.3445, 3.3333, 3.3223, 
    3.3113, 3.3003, 3.2895, 3.2787, 3.268, 3.2573, 3.2468, 3.2362, 3.2258, 
    3.2154, 3.2051, 3.1949, 3.1847, 3.1746, 3.1646, 3.1546, 3.1447, 3.1348, 
    3.125, 3.1153, 3.1056, 3.096, 3.0864, 3.0769, 3.0675, 3.0581, 3.0488, 
    3.0395, 3.0303, 3.0211, 3.012, 3.003, 2.994, 2.9851, 2.9762, 2.9674, 
    2.9586, 2.9499, 2.9412, 2.9326, 2.924, 2.9155, 2.907, 2.8986, 2.8902, 
    2.8818, 2.8736, 2.8653, 2.8571, 2.849, 2.8409, 2.8329, 2.8249, 2.8169, 
    2.809, 2.8011, 2.7933, 2.7855, 2.7778, 2.7701, 2.7624, 2.7548, 2.7473, 
    2.7397, 2.7322, 2.7248, 2.7174, 2.71, 2.7027, 2.6954, 2.6882, 2.681, 
    2.6738, 2.6667, 2.6596, 2.6525, 2.6455, 2.6385, 2.6316, 2.6247, 2.6178, 
    2.611, 2.6042, 2.5974, 2.5907, 2.584, 2.5773, 2.5707, 2.5641, 2.5575, 
    2.551, 2.5445, 2.5381, 2.5316, 2.5253, 2.5189, 2.5126, 2.5063, 2.5, 2.49, 
    2.48, 2.47, 2.46, 2.45, 2.44, 2.43, 2.42, 2.41, 2.4, 2.39, 2.38, 2.37, 
    2.36, 2.35, 2.34, 2.33, 2.32, 2.31, 2.3, 2.29, 2.28, 2.27, 2.26, 2.25, 
    2.24, 2.23, 2.22, 2.21, 2.2, 2.19, 2.18, 2.17, 2.16, 2.15, 2.14, 2.13, 
    2.12, 2.11, 2.1, 2.09, 2.08, 2.07, 2.06, 2.05, 2.04, 2.03, 2.02, 2.01, 2, 
    1.99, 1.98, 1.97, 1.96, 1.95, 1.94, 1.93, 1.92, 1.91, 1.9, 1.89, 1.88, 
    1.87, 1.86, 1.85, 1.84, 1.83, 1.82, 1.81, 1.8, 1.79, 1.78, 1.77, 1.76, 
    1.75, 1.74, 1.73, 1.72, 1.71, 1.7, 1.69, 1.68, 1.67, 1.66, 1.65, 1.64, 
    1.63, 1.62, 1.61, 1.6, 1.59, 1.58, 1.57, 1.56, 1.55, 1.54, 1.53, 1.52, 
    1.51, 1.5, 1.49, 1.48, 1.47, 1.46, 1.45, 1.44, 1.43, 1.42, 1.41, 1.4, 
    1.39, 1.38, 1.37, 1.36, 1.35, 1.34, 1.33, 1.32, 1.31, 1.3, 1.29, 1.28, 
    1.27, 1.26, 1.25, 1.24, 1.23, 1.22, 1.21, 1.2, 1.19, 1.18, 1.17, 1.16, 
    1.15, 1.14, 1.13, 1.12, 1.11, 1.1, 1.09, 1.08, 1.07, 1.06, 1.05, 1.04, 
    1.03, 1.02, 1.01, 1, 0.99, 0.98, 0.97, 0.96, 0.95, 0.94, 0.93, 0.92, 
    0.91, 0.9, 0.89, 0.88, 0.87, 0.86, 0.85, 0.84, 0.83, 0.82, 0.81, 0.8, 
    0.79, 0.78, 0.77, 0.76, 0.75, 0.74, 0.73, 0.72, 0.71, 0.7, 0.69, 0.68, 
    0.67, 0.66, 0.65, 0.64, 0.63, 0.62, 0.61, 0.6, 0.59, 0.58, 0.57, 0.56, 
    0.55, 0.54, 0.53, 0.52, 0.51, 0.5, 0.49, 0.48, 0.47, 0.46, 0.45, 0.44, 
    0.43, 0.42, 0.41, 0.4, 0.39, 0.38, 0.37, 0.36, 0.35, 0.34, 0.33, 0.32, 
    0.31, 0.3, 0.29, 0.28, 0.27, 0.26, 0.25, 0.24, 0.23, 0.22, 0.21 ,
// Copy data from 0.21 um to 0.20 um
	0.20;

 idx_rfr_Fe2O3_eray_roush_rl = 4.916, 5.023, 5.148, 5.292, 5.507, 5.727, 
    6.062, 6.523, 7.11, 7.971, 9.429, 10.555, 7.255, 3.189, 1.513, 0.869, 
    0.706, 0.668, 0.572, 0.489, 0.459, 0.516, 0.599, 0.955, 1.459, 1.862, 
    2.22, 2.513, 2.787, 3.064, 3.336, 3.648, 3.969, 4.568, 4.909, 3.901, 
    2.575, 1.561, 0.989, 0.715, 0.526, 0.42, 0.36, 0.343, 0.329, 0.315, 
    0.319, 0.379, 0.55, 0.787, 0.959, 1.064, 1.182, 1.27, 1.345, 1.407, 
    1.467, 1.522, 1.576, 1.622, 1.665, 1.7, 1.731, 1.765, 1.797, 1.827, 
    1.848, 1.868, 1.89, 1.913, 1.934, 1.948, 1.96, 1.978, 1.994, 2.006, 
    2.018, 2.03, 2.048, 2.064, 2.077, 2.085, 2.095, 2.108, 2.115, 2.124, 
    2.135, 2.146, 2.159, 2.167, 2.174, 2.181, 2.187, 2.193, 2.199, 2.205, 
    2.211, 2.216, 2.221, 2.226, 2.231, 2.236, 2.24, 2.244, 2.249, 2.253, 
    2.257, 2.262, 2.266, 2.269, 2.272, 2.276, 2.28, 2.283, 2.286, 2.29, 
    2.293, 2.296, 2.299, 2.302, 2.305, 2.307, 2.31, 2.312, 2.314, 2.316, 
    2.319, 2.322, 2.324, 2.326, 2.327, 2.329, 2.331, 2.333, 2.334, 2.336, 
    2.337, 2.338, 2.339, 2.341, 2.342, 2.343, 2.344, 2.345, 2.347, 2.348, 
    2.35, 2.351, 2.352, 2.354, 2.355, 2.356, 2.357, 2.358, 2.36, 2.361, 
    2.362, 2.362, 2.363, 2.365, 2.366, 2.367, 2.368, 2.369, 2.37, 2.371, 
    2.371, 2.372, 2.372, 2.373, 2.374, 2.375, 2.376, 2.377, 2.377, 2.377, 
    2.378, 2.378, 2.379, 2.379, 2.379, 2.38, 2.38, 2.38, 2.38, 2.38, 2.381, 
    2.382, 2.382, 2.382, 2.382, 2.383, 2.383, 2.383, 2.383, 2.383, 2.383, 
    2.383, 2.384, 2.384, 2.385, 2.385, 2.385, 2.386, 2.386, 2.386, 2.387, 
    2.387, 2.388, 2.388, 2.389, 2.389, 2.389, 2.389, 2.39, 2.39, 2.39, 2.391, 
    2.391, 2.392, 2.392, 2.393, 2.393, 2.393, 2.393, 2.393, 2.394, 2.394, 
    2.394, 2.395, 2.395, 2.396, 2.396, 2.396, 2.396, 2.395, 2.395, 2.394, 
    2.395, 2.395, 2.395, 2.395, 2.395, 2.396, 2.396, 2.396, 2.396, 2.396, 
    2.396, 2.396, 2.396, 2.397, 2.398, 2.399, 2.399, 2.4, 2.4, 2.4, 2.4, 2.4, 
    2.399, 2.399, 2.399, 2.399, 2.399, 2.399, 2.399, 2.4, 2.401, 2.401, 
    2.401, 2.401, 2.402, 2.403, 2.404, 2.404, 2.405, 2.405, 2.406, 2.406, 
    2.406, 2.406, 2.407, 2.408, 2.41, 2.41, 2.411, 2.411, 2.41, 2.41, 2.41, 
    2.41, 2.41, 2.41, 2.41, 2.411, 2.412, 2.412, 2.413, 2.413, 2.413, 2.412, 
    2.411, 2.411, 2.411, 2.411, 2.411, 2.41, 2.41, 2.41, 2.41, 2.411, 2.411, 
    2.412, 2.413, 2.413, 2.412, 2.412, 2.413, 2.414, 2.415, 2.416, 2.416, 
    2.416, 2.416, 2.416, 2.416, 2.417, 2.418, 2.418, 2.418, 2.418, 2.418, 
    2.418, 2.418, 2.419, 2.419, 2.419, 2.419, 2.419, 2.419, 2.419, 2.419, 
    2.42, 2.42, 2.419, 2.419, 2.418, 2.418, 2.418, 2.419, 2.419, 2.42, 2.42, 
    2.42, 2.42, 2.42, 2.42, 2.421, 2.421, 2.421, 2.421, 2.421, 2.421, 2.421, 
    2.422, 2.423, 2.423, 2.422, 2.422, 2.422, 2.422, 2.422, 2.423, 2.424, 
    2.425, 2.425, 2.425, 2.425, 2.425, 2.426, 2.426, 2.426, 2.427, 2.427, 
    2.428, 2.428, 2.428, 2.428, 2.428, 2.428, 2.428, 2.428, 2.428, 2.428, 
    2.428, 2.428, 2.429, 2.429, 2.429, 2.429, 2.429, 2.429, 2.429, 2.429, 
    2.429, 2.43, 2.43, 2.43, 2.43, 2.43, 2.43, 2.43, 2.43, 2.43, 2.43, 2.43, 
    2.43, 2.43, 2.43, 2.43, 2.431, 2.431, 2.431, 2.432, 2.431, 2.431, 2.432, 
    2.432, 2.432, 2.432, 2.432, 2.432, 2.432, 2.433, 2.433, 2.433, 2.434, 
    2.434, 2.434, 2.434, 2.434, 2.434, 2.433, 2.432, 2.431, 2.431, 2.432, 
    2.433, 2.433, 2.434, 2.435, 2.436, 2.437, 2.438, 2.437, 2.438, 2.438, 
    2.438, 2.438, 2.439, 2.439, 2.44, 2.44, 2.44, 2.441, 2.441, 2.441, 2.441, 
    2.442, 2.442, 2.442, 2.442, 2.443, 2.444, 2.445, 2.446, 2.446, 2.446, 
    2.446, 2.447, 2.448, 2.448, 2.449, 2.449, 2.45, 2.451, 2.452, 2.453, 
    2.453, 2.454, 2.454, 2.455, 2.456, 2.457, 2.458, 2.459, 2.46, 2.461, 
    2.463, 2.463, 2.464, 2.465, 2.466, 2.468, 2.47, 2.471, 2.473, 2.473, 
    2.474, 2.476, 2.477, 2.479, 2.48, 2.482, 2.483, 2.486, 2.488, 2.49, 
    2.491, 2.492, 2.494, 2.496, 2.498, 2.5, 2.502, 2.504, 2.507, 2.51, 2.512, 
    2.515, 2.517, 2.52, 2.522, 2.525, 2.527, 2.529, 2.531, 2.533, 2.535, 
    2.537, 2.541, 2.544, 2.547, 2.549, 2.552, 2.555, 2.559, 2.562, 2.566, 
    2.57, 2.575, 2.582, 2.589, 2.596, 2.604, 2.612, 2.621, 2.631, 2.641, 
    2.652, 2.662, 2.675, 2.688, 2.703, 2.719, 2.736, 2.753, 2.775, 2.8, 2.83, 
    2.862, 2.898, 2.931, 2.956, 2.963, 2.951, 2.927, 2.901, 2.885, 2.881, 
    2.887, 2.893, 2.89, 2.876, 2.858, 2.837, 2.809, 2.766, 2.708, 2.638, 
    2.56, 2.475, 2.387, 2.305, 2.243, 2.211, 2.206, 2.219, 2.218, 2.185, 
    2.134, 2.09, 2.049, 1.992, 1.917, 1.828, 1.733, 1.635, 1.517, 1.349, 1.108,
// Copy data from 0.21 um to 0.20 um
	 1.108;

 idx_rfr_Fe2O3_eray_roush_img = 0.14, 0.157, 0.175, 0.193, 0.218, 0.258, 
    0.294, 0.406, 0.636, 1.037, 2.08, 5.441, 9.384, 8.711, 6.919, 5.566, 
    4.534, 3.852, 3.359, 2.824, 2.315, 1.817, 1.275, 0.743, 0.483, 0.364, 
    0.378, 0.441, 0.429, 0.559, 0.7, 0.857, 1.089, 1.585, 2.831, 4.194, 
    4.452, 4.088, 3.531, 3.059, 2.661, 2.317, 1.99, 1.721, 1.477, 1.242, 
    0.98, 0.69, 0.419, 0.262, 0.256, 0.204, 0.171, 0.152, 0.138, 0.123, 
    0.107, 0.095, 0.084, 0.079, 0.076, 0.074, 0.067, 0.06, 0.058, 0.059, 
    0.061, 0.058, 0.054, 0.051, 0.054, 0.055, 0.049, 0.047, 0.046, 0.045, 
    0.044, 0.037, 0.034, 0.034, 0.035, 0.038, 0.033, 0.035, 0.035, 0.03, 
    0.028, 0.03, 0.031, 0.033, 0.035, 0.036, 0.037, 0.037, 0.038, 0.038, 
    0.039, 0.039, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.042, 0.042, 0.042, 0.042, 
    0.043, 0.044, 0.044, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.046, 
    0.047, 0.047, 0.048, 0.048, 0.048, 0.049, 0.049, 0.05, 0.05, 0.05, 0.051, 
    0.051, 0.051, 0.05, 0.051, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.051, 0.051, 0.051, 0.05, 0.051, 0.051, 
    0.051, 0.051, 0.052, 0.052, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.054, 0.054, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.056, 0.056, 0.056, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.054, 0.054, 0.054, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.052, 0.052, 0.052, 0.051, 0.051, 0.051, 0.051, 
    0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.049, 0.05, 0.05, 0.051, 
    0.051, 0.051, 0.051, 0.05, 0.049, 0.049, 0.049, 0.049, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.047, 0.047, 0.046, 0.045, 0.045, 0.044, 0.044, 
    0.045, 0.045, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.045, 0.045, 
    0.044, 0.043, 0.042, 0.042, 0.041, 0.041, 0.041, 0.04, 0.04, 0.039, 
    0.039, 0.04, 0.039, 0.039, 0.039, 0.04, 0.04, 0.039, 0.039, 0.038, 0.039, 
    0.039, 0.04, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.04, 0.04, 0.04, 0.041, 0.042, 0.043, 0.043, 0.043, 0.043, 0.042, 0.042, 
    0.042, 0.042, 0.041, 0.041, 0.04, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.038, 0.037, 0.037, 0.037, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.04, 0.04, 0.04, 0.04, 0.041, 0.041, 0.041, 
    0.04, 0.04, 0.039, 0.038, 0.038, 0.038, 0.039, 0.039, 0.039, 0.039, 
    0.038, 0.038, 0.039, 0.039, 0.039, 0.038, 0.038, 0.037, 0.037, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.037, 0.036, 0.036, 0.037, 0.037, 
    0.037, 0.037, 0.037, 0.037, 0.038, 0.037, 0.038, 0.038, 0.039, 0.039, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.041, 0.04, 0.04, 0.04, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.041, 0.041, 0.041, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.041, 0.041, 0.041, 0.041, 0.041, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.043, 0.043, 0.043, 0.042, 0.04, 0.039, 
    0.038, 0.038, 0.038, 0.037, 0.037, 0.037, 0.038, 0.039, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.037, 0.036, 0.036, 0.036, 0.036, 0.037, 
    0.037, 0.036, 0.036, 0.036, 0.035, 0.035, 0.035, 0.035, 0.034, 0.034, 
    0.035, 0.035, 0.035, 0.034, 0.034, 0.034, 0.033, 0.033, 0.033, 0.033, 
    0.033, 0.033, 0.033, 0.033, 0.033, 0.032, 0.032, 0.032, 0.033, 0.033, 
    0.033, 0.034, 0.033, 0.034, 0.034, 0.034, 0.033, 0.033, 0.034, 0.034, 
    0.035, 0.036, 0.036, 0.036, 0.036, 0.037, 0.037, 0.038, 0.038, 0.039, 
    0.039, 0.04, 0.042, 0.042, 0.043, 0.045, 0.046, 0.048, 0.049, 0.051, 
    0.051, 0.052, 0.053, 0.053, 0.054, 0.056, 0.057, 0.058, 0.058, 0.059, 
    0.059, 0.059, 0.058, 0.057, 0.057, 0.057, 0.058, 0.059, 0.06, 0.061, 
    0.063, 0.066, 0.068, 0.072, 0.075, 0.078, 0.083, 0.089, 0.096, 0.103, 
    0.11, 0.119, 0.134, 0.156, 0.186, 0.229, 0.286, 0.351, 0.413, 0.46, 
    0.492, 0.512, 0.532, 0.56, 0.602, 0.654, 0.707, 0.758, 0.813, 0.873, 
    0.936, 0.993, 1.04, 1.075, 1.096, 1.097, 1.075, 1.034, 0.987, 0.951, 
    0.947, 0.979, 1.018, 1.041, 1.053, 1.076, 1.107, 1.133, 1.148, 1.149, 
    1.145, 1.145, 1.127, 1.048 ,
// Copy data from 0.21 um to 0.20 um
	 1.048 ;

 idx_rfr_Fe2O3_eray_roush_rl_ee = 0.118, 0.124, 0.13, 0.138, 0.15, 0.163, 
    0.183, 0.214, 0.257, 0.328, 0.473, 0.648, 0.668, 0.638, 0.39, 0.248, 
    0.179, 0.146, 0.119, 0.093, 0.076, 0.068, 0.06, 0.051, 0.028, 0.022, 
    0.027, 0.035, 0.041, 0.053, 0.065, 0.081, 0.1, 0.142, 0.21, 0.241, 0.277, 
    0.221, 0.159, 0.12, 0.092, 0.073, 0.059, 0.052, 0.046, 0.04, 0.035, 
    0.032, 0.03, 0.025, 0.022, 0.014, 0.009, 0.008, 0.007, 0.007, 0.007, 
    0.008, 0.008, 0.009, 0.01, 0.01, 0.011, 0.011, 0.012, 0.012, 0.013, 
    0.013, 0.013, 0.014, 0.014, 0.014, 0.015, 0.015, 0.015, 0.016, 0.016, 
    0.016, 0.016, 0.017, 0.017, 0.017, 0.017, 0.018, 0.018, 0.018, 0.018, 
    0.018, 0.019, 0.019, 0.019, 0.019, 0.019, 0.019, 0.02, 0.02, 0.02, 0.02, 
    0.02, 0.02, 0.02, 0.02, 0.021, 0.021, 0.021, 0.021, 0.021, 0.021, 0.021, 
    0.021, 0.021, 0.021, 0.021, 0.022, 0.022, 0.022, 0.022, 0.022, 0.022, 
    0.022, 0.022, 0.022, 0.022, 0.022, 0.022, 0.022, 0.022, 0.022, 0.023, 
    0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 
    0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 
    0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.026, 0.026, 0.026, 0.026, 0.026, 
    0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 
    0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 
    0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.027, 
    0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 
    0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.028, 0.028, 0.028, 0.028, 
    0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 
    0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.03, 0.03, 0.03, 0.03, 0.031, 
    0.031, 0.031, 0.032, 0.032, 0.032, 0.033, 0.033, 0.034, 0.035, 0.035, 
    0.036, 0.038, 0.039, 0.041, 0.042, 0.044, 0.045, 0.046, 0.046, 0.046, 
    0.047, 0.048, 0.05, 0.052, 0.054, 0.056, 0.058, 0.06, 0.063, 0.065, 
    0.067, 0.068, 0.068, 0.067, 0.065, 0.062, 0.059, 0.057, 0.057, 0.059, 
    0.061, 0.062, 0.063, 0.064, 0.066, 0.067, 0.068, 0.067, 0.067, 0.066, 
    0.069, 0.066 ,
// Copy data from 0.21 um to 0.20 um
	0.066 ;	

 idx_rfr_Fe2O3_eray_roush_img_ee = 0.014, 0.016, 0.018, 0.021, 0.024, 0.029, 
    0.034, 0.048, 0.079, 0.137, 0.3, 0.752, 0.823, 0.641, 0.446, 0.337, 0.27, 
    0.228, 0.199, 0.168, 0.14, 0.112, 0.08, 0.029, 0.022, 0.024, 0.027, 
    0.033, 0.034, 0.045, 0.057, 0.072, 0.093, 0.139, 0.214, 0.19, 0.244, 
    0.237, 0.207, 0.18, 0.159, 0.141, 0.124, 0.111, 0.1, 0.09, 0.079, 0.068, 
    0.052, 0.027, 0.009, 0.005, 0.009, 0.009, 0.009, 0.008, 0.007, 0.006, 
    0.006, 0.005, 0.005, 0.005, 0.005, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.002, 0.003, 0.003, 0.003, 0.002, 0.003, 0.003, 0.002, 0.002, 0.002, 
    0.002, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.003, 0.003, 0.003, 0.003, 0.003, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.002, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.005, 0.005, 0.005, 0.005, 
    0.005, 0.005, 0.005, 0.005, 0.004, 0.005, 0.005, 0.005, 0.005, 0.005, 
    0.005, 0.005, 0.005, 0.006, 0.006, 0.006, 0.007, 0.007, 0.008, 0.008, 
    0.009, 0.01, 0.011, 0.013, 0.015, 0.019, 0.023, 0.029, 0.033, 0.037, 
    0.039, 0.04, 0.042, 0.044, 0.046, 0.05, 0.053, 0.056, 0.059, 0.061, 
    0.064, 0.065, 0.065, 0.064, 0.062, 0.06, 0.057, 0.054, 0.052, 0.051, 
    0.051, 0.052, 0.052, 0.05, 0.049, 0.047, 0.045, 0.041, 0.037, 0.031, 
    0.025, 0.018, 0.025, 0.035 ,
// Copy data from 0.21 um to 0.20 um
	0.035 ;

 idx_rfr_Fe2O3_eray_roush_nr = 0.44077, 0.44879, 0.45795, 0.4681, 0.48255, 
    0.49675, 0.5168, 0.54245, 0.5723, 0.611, 0.66825, 0.7426, 0.8153, 0.8643, 
    0.889, 0.89975, 0.88045, 0.8492, 0.83465, 0.80945, 0.7563, 0.6336, 
    0.43055, 0.1289, 0.07185, 0.10655, 0.157, 0.20005, 0.2346, 0.27395, 
    0.31055, 0.34905, 0.3888, 0.4571, 0.54475, 0.6269, 0.6858, 0.73315, 
    0.7605, 0.76895, 0.77785, 0.7741, 0.75355, 0.714, 0.6691, 0.61785, 
    0.53115, 0.3679, 0.151, 0.036, 0.0177, 0.0109, 0.0133, 0.0189, 0.02555, 
    0.0317, 0.03825, 0.0449, 0.0518, 0.0581, 0.06395, 0.06895, 0.0733, 
    0.07805, 0.08275, 0.08715, 0.09035, 0.0932, 0.0964, 0.0999, 0.103, 
    0.10505, 0.10685, 0.10955, 0.11185, 0.1137, 0.1155, 0.1172, 0.1198, 
    0.12225, 0.1242, 0.1253, 0.12685, 0.1287, 0.12975, 0.13115, 0.1328, 
    0.13435, 0.1363, 0.13745, 0.1385, 0.13955, 0.14045, 0.14135, 0.1423, 
    0.1432, 0.144, 0.14475, 0.1455, 0.14625, 0.14695, 0.14765, 0.1483, 
    0.1489, 0.14955, 0.15025, 0.15085, 0.15145, 0.15205, 0.15255, 0.15305, 
    0.1536, 0.1541, 0.1546, 0.1551, 0.1556, 0.15605, 0.15655, 0.157, 0.1574, 
    0.1578, 0.15815, 0.1585, 0.1588, 0.1591, 0.15945, 0.15985, 0.16025, 
    0.16055, 0.16085, 0.1611, 0.16135, 0.16165, 0.1619, 0.1621, 0.16235, 
    0.16255, 0.1627, 0.16285, 0.16305, 0.1632, 0.1634, 0.16355, 0.1637, 
    0.1639, 0.16405, 0.1643, 0.1645, 0.1647, 0.1649, 0.16505, 0.16525, 
    0.16545, 0.1656, 0.1658, 0.1659, 0.16605, 0.16615, 0.1663, 0.1665, 
    0.16665, 0.1668, 0.167, 0.16715, 0.1673, 0.16735, 0.1674, 0.1675, 0.1676, 
    0.16775, 0.16785, 0.16795, 0.1681, 0.16825, 0.1683, 0.16835, 0.1684, 
    0.16845, 0.16855, 0.1686, 0.16865, 0.1687, 0.1687, 0.1687, 0.1687, 
    0.1688, 0.1689, 0.16895, 0.169, 0.16905, 0.16905, 0.1691, 0.1691, 0.1691, 
    0.1691, 0.16915, 0.1692, 0.1692, 0.16925, 0.16935, 0.1694, 0.1694, 
    0.16945, 0.1695, 0.16955, 0.1696, 0.16965, 0.16975, 0.1698, 0.1699, 
    0.16995, 0.17, 0.17005, 0.17005, 0.1701, 0.17015, 0.1702, 0.17025, 
    0.1703, 0.1704, 0.17045, 0.1705, 0.17055, 0.1706, 0.1706, 0.1706, 
    0.17065, 0.1707, 0.17075, 0.1708, 0.17085, 0.17095, 0.171, 0.17105, 
    0.171, 0.1709, 0.1708, 0.17075, 0.1708, 0.17085, 0.17085, 0.17085, 
    0.1709, 0.17095, 0.17095, 0.17095, 0.17095, 0.17095, 0.17095, 0.17095, 
    0.171, 0.1711, 0.17125, 0.1714, 0.17145, 0.17155, 0.17155, 0.1715, 
    0.1715, 0.1715, 0.17145, 0.17145, 0.1714, 0.1714, 0.17135, 0.17135, 
    0.1714, 0.1715, 0.1716, 0.17165, 0.17165, 0.1717, 0.1718, 0.17195, 
    0.17205, 0.1721, 0.17215, 0.17225, 0.17235, 0.1724, 0.1724, 0.1724, 
    0.17255, 0.1727, 0.17285, 0.1729, 0.173, 0.173, 0.17295, 0.17295, 0.173, 
    0.173, 0.17295, 0.17295, 0.17295, 0.17305, 0.17315, 0.17325, 0.1733, 
    0.1734, 0.1734, 0.17325, 0.17315, 0.1731, 0.17305, 0.17305, 0.17305, 
    0.173, 0.173, 0.17295, 0.17295, 0.173, 0.1731, 0.17325, 0.17335, 0.1733, 
    0.17325, 0.17325, 0.17335, 0.1735, 0.1736, 0.1737, 0.1737, 0.17375, 
    0.17375, 0.1737, 0.1738, 0.1739, 0.174, 0.17405, 0.1741, 0.1741, 0.17405, 
    0.17405, 0.1741, 0.17415, 0.17415, 0.17415, 0.1742, 0.1742, 0.17425, 
    0.17425, 0.17425, 0.1743, 0.1743, 0.1742, 0.17415, 0.1741, 0.17405, 
    0.17405, 0.17415, 0.17425, 0.17435, 0.1744, 0.1744, 0.17435, 0.17435, 
    0.1744, 0.17445, 0.1745, 0.1745, 0.17445, 0.17445, 0.17445, 0.1745, 
    0.17465, 0.17475, 0.1747, 0.17465, 0.17465, 0.17465, 0.17465, 0.17465, 
    0.1748, 0.17495, 0.17505, 0.175, 0.175, 0.17505, 0.1751, 0.17515, 0.1752, 
    0.1752, 0.1753, 0.1754, 0.17545, 0.1755, 0.1755, 0.17545, 0.17545, 
    0.17545, 0.1755, 0.1755, 0.1755, 0.1755, 0.1755, 0.17555, 0.1756, 0.1756, 
    0.1756, 0.1756, 0.17565, 0.1757, 0.1757, 0.1757, 0.1757, 0.17575, 
    0.17575, 0.17575, 0.17575, 0.1758, 0.1758, 0.1758, 0.1758, 0.1758, 
    0.1758, 0.1758, 0.1758, 0.17585, 0.17585, 0.17585, 0.1759, 0.1759, 
    0.17595, 0.176, 0.176, 0.176, 0.176, 0.17605, 0.17605, 0.17605, 0.17605, 
    0.1761, 0.1761, 0.17615, 0.1762, 0.17625, 0.1763, 0.1763, 0.1763, 0.1763, 
    0.1763, 0.1763, 0.1762, 0.17605, 0.17595, 0.1759, 0.17605, 0.17615, 
    0.17625, 0.17635, 0.1765, 0.17665, 0.1768, 0.17685, 0.1768, 0.17685, 
    0.1769, 0.1769, 0.17695, 0.177, 0.17705, 0.17715, 0.1772, 0.17725, 
    0.1773, 0.17735, 0.1774, 0.1774, 0.17745, 0.17745, 0.17745, 0.1775, 
    0.1776, 0.1777, 0.17785, 0.178, 0.178, 0.178, 0.17805, 0.17815, 0.17825, 
    0.1783, 0.1784, 0.1785, 0.1786, 0.17875, 0.17885, 0.179, 0.17905, 0.1791, 
    0.1792, 0.1793, 0.1794, 0.17955, 0.1797, 0.1799, 0.18005, 0.1802, 0.1804, 
    0.18045, 0.1806, 0.1807, 0.1809, 0.1811, 0.18135, 0.18155, 0.1818, 
    0.1819, 0.18205, 0.18225, 0.18245, 0.18265, 0.18285, 0.18305, 0.1833, 
    0.18365, 0.18395, 0.1842, 0.1844, 0.18455, 0.1848, 0.18505, 0.18535, 
    0.1857, 0.186, 0.1863, 0.18665, 0.18705, 0.1874, 0.18775, 0.18805, 
    0.18845, 0.18885, 0.1892, 0.18955, 0.1898, 0.19005, 0.19035, 0.19065, 
    0.191, 0.19145, 0.1919, 0.1923, 0.1927, 0.1931, 0.1935, 0.194, 0.19445, 
    0.195, 0.19555, 0.19625, 0.19715, 0.19815, 0.1992, 0.20025, 0.2014, 
    0.20265, 0.204, 0.2054, 0.20685, 0.20835, 0.21005, 0.2119, 0.2139, 
    0.21615, 0.21845, 0.22085, 0.22375, 0.2272, 0.23135, 0.23585, 0.2409, 
    0.24605, 0.25055, 0.25345, 0.2542, 0.2532, 0.2516, 0.2506, 0.25115, 
    0.2534, 0.25645, 0.2592, 0.2611, 0.26265, 0.26455, 0.2664, 0.2675, 
    0.2671, 0.2652, 0.26175, 0.25655, 0.24895, 0.23885, 0.22775, 0.2183, 
    0.21305, 0.2137, 0.2179, 0.22035, 0.2194, 0.2177, 0.2181, 0.21925, 
    0.2192, 0.2173, 0.21345, 0.2098, 0.2086, 0.20735, 0.20265 ,
// Copy data from 0.21 um to 0.20 um
	0.20265 ;

 bnd_wvn_Fe2O3_oray_roush = 180, 190, 200, 210, 220, 230, 240, 250, 260, 270, 
    280, 290, 300, 310, 320, 330, 340, 350, 360, 370, 380, 390, 400, 410, 
    420, 430, 440, 450, 460, 470, 480, 490, 500, 510, 520, 530, 540, 550, 
    560, 570, 580, 590, 600, 610, 620, 630, 640, 650, 660, 670, 680, 690, 
    700, 710, 720, 730, 740, 750, 760, 770, 780, 790, 800, 810, 820, 830, 
    840, 850, 860, 870, 880, 890, 900, 910, 920, 930, 940, 950, 960, 970, 
    980, 990, 1000, 1010, 1020, 1030, 1040, 1050, 1060, 1070, 1080, 1090, 
    1100, 1110, 1120, 1130, 1140, 1150, 1160, 1170, 1180, 1190, 1200, 1210, 
    1220, 1230, 1240, 1250, 1260, 1270, 1280, 1290, 1300, 1310, 1320, 1330, 
    1340, 1350, 1360, 1370, 1380, 1390, 1400, 1410, 1420, 1430, 1440, 1450, 
    1460, 1470, 1480, 1490, 1500, 1510, 1520, 1530, 1540, 1550, 1560, 1570, 
    1580, 1590, 1600, 1610, 1620, 1630, 1640, 1650, 1660, 1670, 1680, 1690, 
    1700, 1710, 1720, 1730, 1740, 1750, 1760, 1770, 1780, 1790, 1800, 1810, 
    1820, 1830, 1840, 1850, 1860, 1870, 1880, 1890, 1900, 1910, 1920, 1930, 
    1940, 1950, 1960, 1970, 1980, 1990, 2000, 2010, 2020, 2030, 2040, 2050, 
    2060, 2070, 2080, 2090, 2100, 2110, 2120, 2130, 2140, 2150, 2160, 2170, 
    2180, 2190, 2200, 2210, 2220, 2230, 2240, 2250, 2260, 2270, 2280, 2290, 
    2300, 2310, 2320, 2330, 2340, 2350, 2360, 2370, 2380, 2390, 2400, 2410, 
    2420, 2430, 2440, 2450, 2460, 2470, 2480, 2490, 2500, 2510, 2520, 2530, 
    2540, 2550, 2560, 2570, 2580, 2590, 2600, 2610, 2620, 2630, 2640, 2650, 
    2660, 2670, 2680, 2690, 2700, 2710, 2720, 2730, 2740, 2750, 2760, 2770, 
    2780, 2790, 2800, 2810, 2820, 2830, 2840, 2850, 2860, 2870, 2880, 2890, 
    2900, 2910, 2920, 2930, 2940, 2950, 2960, 2970, 2980, 2990, 3000, 3010, 
    3020, 3030, 3040, 3050, 3060, 3070, 3080, 3090, 3100, 3110, 3120, 3130, 
    3140, 3150, 3160, 3170, 3180, 3190, 3200, 3210, 3220, 3230, 3240, 3250, 
    3260, 3270, 3280, 3290, 3300, 3310, 3320, 3330, 3340, 3350, 3360, 3370, 
    3380, 3390, 3400, 3410, 3420, 3430, 3440, 3450, 3460, 3470, 3480, 3490, 
    3500, 3510, 3520, 3530, 3540, 3550, 3560, 3570, 3580, 3590, 3600, 3610, 
    3620, 3630, 3640, 3650, 3660, 3670, 3680, 3690, 3700, 3710, 3720, 3730, 
    3740, 3750, 3760, 3770, 3780, 3790, 3800, 3810, 3820, 3830, 3840, 3850, 
    3860, 3870, 3880, 3890, 3900, 3910, 3920, 3930, 3940, 3950, 3960, 3970, 
    3980, 3990, 4000, 4016.06, 4032.26, 4048.58, 4065.04, 4081.63, 4098.36, 
    4115.23, 4132.23, 4149.38, 4166.67, 4184.1, 4201.68, 4219.41, 4237.29, 
    4255.32, 4273.5, 4291.85, 4310.34, 4329, 4347.83, 4366.81, 4385.96, 
    4405.29, 4424.78, 4444.44, 4464.29, 4484.3, 4504.5, 4524.89, 4545.45, 
    4566.21, 4587.16, 4608.29, 4629.63, 4651.16, 4672.9, 4694.84, 4716.98, 
    4739.34, 4761.9, 4784.69, 4807.69, 4830.92, 4854.37, 4878.05, 4901.96, 
    4926.11, 4950.5, 4975.12, 5000, 5025.13, 5050.51, 5076.14, 5102.04, 
    5128.21, 5154.64, 5181.35, 5208.33, 5235.6, 5263.16, 5291.01, 5319.15, 
    5347.59, 5376.34, 5405.41, 5434.78, 5464.48, 5494.51, 5524.86, 5555.56, 
    5586.59, 5617.98, 5649.72, 5681.82, 5714.29, 5747.13, 5780.35, 5813.95, 
    5847.95, 5882.35, 5917.16, 5952.38, 5988.02, 6024.1, 6060.61, 6097.56, 
    6134.97, 6172.84, 6211.18, 6250, 6289.31, 6329.11, 6369.43, 6410.26, 
    6451.61, 6493.51, 6535.95, 6578.95, 6622.52, 6666.67, 6711.41, 6756.76, 
    6802.72, 6849.32, 6896.55, 6944.44, 6993.01, 7042.25, 7092.2, 7142.86, 
    7194.24, 7246.38, 7299.27, 7352.94, 7407.41, 7462.69, 7518.8, 7575.76, 
    7633.59, 7692.31, 7751.94, 7812.5, 7874.02, 7936.51, 8000, 8064.52, 
    8130.08, 8196.72, 8264.46, 8333.33, 8403.36, 8474.58, 8547.01, 8620.69, 
    8695.65, 8771.93, 8849.56, 8928.57, 9009.01, 9090.91, 9174.31, 9259.26, 
    9345.79, 9433.96, 9523.81, 9615.38, 9708.74, 9803.92, 9900.99, 10000, 
    10101.01, 10204.08, 10309.28, 10416.67, 10526.32, 10638.3, 10752.69, 
    10869.57, 10989.01, 11111.11, 11235.96, 11363.64, 11494.25, 11627.91, 
    11764.71, 11904.76, 12048.19, 12195.12, 12345.68, 12500, 12658.23, 
    12820.51, 12987.01, 13157.89, 13333.33, 13513.51, 13698.63, 13888.89, 
    14084.51, 14285.71, 14492.75, 14705.88, 14925.37, 15151.52, 15384.62, 
    15625, 15873.02, 16129.03, 16393.44, 16666.67, 16949.15, 17241.38, 
    17543.86, 17857.14, 18181.82, 18518.52, 18867.92, 19230.77, 19607.84, 
    20000, 20408.16, 20833.33, 21276.6, 21739.13, 22222.22, 22727.27, 
    23255.81, 23809.52, 24390.24, 25000, 25641.03, 26315.79, 27027.03, 
    27777.78, 28571.43, 29411.76, 30303.03, 31250, 32258.06, 33333.33, 
    34482.76, 35714.29, 37037.04, 38461.54, 40000, 41666.67, 43478.26, 
    45454.55, 47619.05, 50000 ;

 idx_rfr_Fe2O3_oray_roush_rl = 5.658, 5.844, 6.094, 6.359, 6.789, 7.022, 
    6.649, 7.29, 8.312, 9.433, 11.932, 12.585, 6.494, 2.681, 1.402, 1.005, 
    0.846, 0.808, 1.03, 1.554, 2.383, 3.262, 4.1, 4.966, 6.229, 7.431, 4.992, 
    2.23, 1.268, 1.015, 0.902, 1.105, 1.764, 2.673, 2.82, 2.007, 1.265, 
    0.787, 0.522, 0.395, 0.342, 0.318, 0.304, 0.307, 0.327, 0.361, 0.403, 
    0.478, 0.601, 0.754, 0.91, 1.037, 1.145, 1.238, 1.322, 1.399, 1.471, 
    1.536, 1.597, 1.653, 1.702, 1.745, 1.786, 1.823, 1.857, 1.891, 1.921, 
    1.949, 1.974, 1.999, 2.023, 2.045, 2.065, 2.081, 2.095, 2.11, 2.126, 
    2.141, 2.155, 2.17, 2.185, 2.199, 2.212, 2.224, 2.236, 2.246, 2.256, 
    2.265, 2.275, 2.284, 2.294, 2.303, 2.312, 2.321, 2.329, 2.337, 2.344, 
    2.349, 2.356, 2.363, 2.369, 2.375, 2.381, 2.386, 2.392, 2.398, 2.404, 
    2.409, 2.414, 2.418, 2.423, 2.428, 2.433, 2.438, 2.443, 2.447, 2.452, 
    2.457, 2.462, 2.466, 2.469, 2.474, 2.477, 2.481, 2.485, 2.488, 2.491, 
    2.494, 2.498, 2.5, 2.503, 2.505, 2.508, 2.511, 2.514, 2.516, 2.517, 2.52, 
    2.522, 2.524, 2.525, 2.527, 2.529, 2.532, 2.534, 2.536, 2.539, 2.541, 
    2.542, 2.543, 2.545, 2.547, 2.549, 2.551, 2.552, 2.554, 2.556, 2.557, 
    2.559, 2.56, 2.561, 2.562, 2.564, 2.565, 2.567, 2.568, 2.569, 2.57, 
    2.572, 2.573, 2.575, 2.575, 2.576, 2.578, 2.579, 2.58, 2.581, 2.582, 
    2.583, 2.584, 2.585, 2.586, 2.587, 2.588, 2.588, 2.59, 2.591, 2.592, 
    2.593, 2.593, 2.595, 2.595, 2.596, 2.597, 2.598, 2.598, 2.599, 2.6, 
    2.601, 2.602, 2.602, 2.603, 2.604, 2.604, 2.605, 2.605, 2.606, 2.607, 
    2.607, 2.608, 2.609, 2.609, 2.61, 2.611, 2.612, 2.613, 2.615, 2.615, 
    2.616, 2.616, 2.615, 2.615, 2.616, 2.618, 2.619, 2.619, 2.62, 2.62, 
    2.621, 2.622, 2.623, 2.623, 2.624, 2.624, 2.624, 2.625, 2.625, 2.625, 
    2.626, 2.627, 2.627, 2.627, 2.628, 2.628, 2.628, 2.629, 2.63, 2.63, 
    2.631, 2.631, 2.631, 2.632, 2.632, 2.633, 2.633, 2.634, 2.634, 2.634, 
    2.635, 2.635, 2.635, 2.635, 2.635, 2.636, 2.637, 2.637, 2.638, 2.638, 
    2.638, 2.639, 2.639, 2.639, 2.64, 2.64, 2.64, 2.641, 2.64, 2.641, 2.641, 
    2.641, 2.641, 2.641, 2.641, 2.64, 2.64, 2.642, 2.642, 2.642, 2.642, 
    2.643, 2.643, 2.643, 2.643, 2.643, 2.644, 2.644, 2.644, 2.644, 2.645, 
    2.645, 2.646, 2.646, 2.646, 2.646, 2.647, 2.647, 2.648, 2.648, 2.648, 
    2.648, 2.648, 2.648, 2.649, 2.649, 2.65, 2.65, 2.65, 2.65, 2.65, 2.65, 
    2.65, 2.65, 2.65, 2.65, 2.65, 2.651, 2.651, 2.651, 2.652, 2.652, 2.652, 
    2.652, 2.653, 2.653, 2.653, 2.653, 2.654, 2.654, 2.654, 2.655, 2.655, 
    2.655, 2.655, 2.656, 2.656, 2.655, 2.655, 2.656, 2.656, 2.657, 2.657, 
    2.657, 2.657, 2.657, 2.657, 2.658, 2.659, 2.659, 2.658, 2.657, 2.657, 
    2.658, 2.659, 2.659, 2.659, 2.659, 2.659, 2.659, 2.659, 2.659, 2.659, 
    2.659, 2.658, 2.658, 2.658, 2.658, 2.658, 2.657, 2.657, 2.657, 2.658, 
    2.658, 2.658, 2.658, 2.659, 2.659, 2.66, 2.66, 2.659, 2.659, 2.659, 2.66, 
    2.66, 2.66, 2.66, 2.66, 2.661, 2.661, 2.661, 2.661, 2.661, 2.661, 2.662, 
    2.662, 2.662, 2.662, 2.662, 2.662, 2.662, 2.662, 2.662, 2.662, 2.662, 
    2.662, 2.663, 2.663, 2.663, 2.663, 2.663, 2.663, 2.663, 2.664, 2.664, 
    2.664, 2.664, 2.664, 2.664, 2.664, 2.665, 2.665, 2.665, 2.665, 2.665, 
    2.665, 2.666, 2.666, 2.667, 2.667, 2.667, 2.667, 2.667, 2.667, 2.667, 
    2.666, 2.665, 2.664, 2.664, 2.665, 2.666, 2.667, 2.668, 2.669, 2.67, 
    2.671, 2.672, 2.671, 2.672, 2.672, 2.673, 2.673, 2.673, 2.674, 2.674, 
    2.675, 2.676, 2.676, 2.676, 2.677, 2.677, 2.677, 2.677, 2.677, 2.678, 
    2.679, 2.68, 2.681, 2.682, 2.682, 2.682, 2.683, 2.683, 2.684, 2.685, 
    2.686, 2.686, 2.687, 2.689, 2.69, 2.691, 2.692, 2.692, 2.693, 2.693, 
    2.695, 2.696, 2.697, 2.699, 2.7, 2.702, 2.703, 2.704, 2.705, 2.706, 
    2.708, 2.709, 2.712, 2.714, 2.715, 2.716, 2.718, 2.719, 2.721, 2.723, 
    2.725, 2.727, 2.729, 2.732, 2.734, 2.737, 2.739, 2.74, 2.742, 2.745, 
    2.747, 2.75, 2.753, 2.755, 2.759, 2.762, 2.765, 2.768, 2.771, 2.775, 
    2.778, 2.781, 2.784, 2.787, 2.789, 2.791, 2.794, 2.798, 2.801, 2.805, 
    2.809, 2.813, 2.816, 2.82, 2.824, 2.828, 2.833, 2.838, 2.845, 2.853, 
    2.862, 2.872, 2.882, 2.892, 2.903, 2.916, 2.929, 2.942, 2.956, 2.972, 
    2.99, 3.008, 3.029, 3.051, 3.074, 3.102, 3.135, 3.175, 3.218, 3.265, 
    3.312, 3.348, 3.361, 3.348, 3.318, 3.286, 3.266, 3.262, 3.272, 3.282, 
    3.28, 3.264, 3.242, 3.217, 3.181, 3.126, 3.052, 2.962, 2.863, 2.756, 
    2.645, 2.545, 2.47, 2.433, 2.43, 2.45, 2.454, 2.416, 2.357, 2.307, 2.261, 
    2.197, 2.11, 2.007, 1.899, 1.79, 1.659, 1.471, 1.202, 1.202 ;

 idx_rfr_Fe2O3_oray_roush_img =
// csz++
// As supplied by Roush, the first four values had negative refractive indices
// Replace with absoluted values of same to prevent problems downstream
//	 -0.144, -0.148, -0.117, -0.074, 0.03, 0.668, 
    +0.144, +0.148, +0.117, +0.074, 0.03, 0.668, 
    0.601, 0.132, 0.389, 0.782, 2.15, 8.306, 11.145, 9.062, 6.922, 5.382, 
    4.284, 3.245, 2.254, 1.39, 0.803, 0.656, 0.718, 0.982, 1.587, 4.077, 
    6.991, 6.303, 4.993, 4.068, 3.328, 2.553, 2.054, 2.292, 3.368, 3.911, 
    3.791, 3.436, 3.035, 2.669, 2.358, 2.096, 1.855, 1.624, 1.406, 1.201, 
    0.994, 0.779, 0.586, 0.44, 0.35, 0.297, 0.256, 0.221, 0.192, 0.167, 
    0.147, 0.132, 0.119, 0.111, 0.106, 0.102, 0.097, 0.093, 0.088, 0.085, 
    0.083, 0.081, 0.08, 0.077, 0.076, 0.077, 0.078, 0.079, 0.076, 0.072, 
    0.069, 0.066, 0.064, 0.06, 0.058, 0.057, 0.056, 0.055, 0.055, 0.055, 
    0.054, 0.052, 0.05, 0.048, 0.047, 0.046, 0.045, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.043, 0.042, 0.041, 0.04, 0.039, 0.039, 0.038, 0.037, 
    0.036, 0.036, 0.035, 0.035, 0.034, 0.033, 0.032, 0.031, 0.031, 0.031, 
    0.03, 0.029, 0.029, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.031, 0.031, 
    0.031, 0.032, 0.032, 0.032, 0.032, 0.031, 0.032, 0.033, 0.033, 0.033, 
    0.033, 0.033, 0.033, 0.033, 0.032, 0.032, 0.031, 0.031, 0.031, 0.032, 
    0.032, 0.032, 0.032, 0.031, 0.031, 0.032, 0.032, 0.032, 0.031, 0.032, 
    0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.03, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.029, 0.029, 
    0.029, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.029, 0.03, 0.03, 0.03, 
    0.029, 0.028, 0.028, 0.028, 0.029, 0.029, 0.028, 0.028, 0.029, 0.029, 
    0.029, 0.029, 0.029, 0.029, 0.029, 0.03, 0.03, 0.029, 0.03, 0.029, 0.03, 
    0.03, 0.03, 0.029, 0.029, 0.029, 0.029, 0.03, 0.03, 0.03, 0.03, 0.029, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.031, 0.031, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.031, 0.031, 0.031, 0.031, 0.031, 0.032, 
    0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.032, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.03, 0.03, 0.03, 0.031, 
    0.031, 0.031, 0.031, 0.032, 0.031, 0.031, 0.031, 0.031, 0.032, 0.032, 
    0.032, 0.032, 0.032, 0.032, 0.032, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.032, 0.032, 0.032, 0.032, 
    0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.033, 
    0.034, 0.034, 0.034, 0.033, 0.033, 0.033, 0.034, 0.034, 0.034, 0.035, 
    0.035, 0.035, 0.035, 0.035, 0.036, 0.036, 0.036, 0.035, 0.036, 0.036, 
    0.035, 0.035, 0.034, 0.034, 0.034, 0.034, 0.033, 0.034, 0.034, 0.034, 
    0.035, 0.035, 0.035, 0.034, 0.034, 0.034, 0.035, 0.034, 0.034, 0.034, 
    0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 
    0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 
    0.033, 0.033, 0.033, 0.033, 0.033, 0.032, 0.033, 0.033, 0.033, 0.033, 
    0.032, 0.032, 0.032, 0.032, 0.032, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.031, 0.029, 
    0.027, 0.026, 0.026, 0.025, 0.025, 0.024, 0.025, 0.026, 0.026, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.023, 0.023, 0.022, 0.021, 0.02, 0.02, 0.02, 0.021, 
    0.021, 0.02, 0.019, 0.019, 0.019, 0.018, 0.018, 0.017, 0.017, 0.017, 
    0.017, 0.017, 0.017, 0.016, 0.015, 0.015, 0.014, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.012, 0.011, 0.01, 0.01, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.01, 0.01, 0.009, 0.009, 0.01, 0.01, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.012, 
    0.013, 0.014, 0.015, 0.015, 0.017, 0.018, 0.02, 0.021, 0.022, 0.023, 
    0.023, 0.023, 0.024, 0.024, 0.026, 0.026, 0.026, 0.027, 0.027, 0.026, 
    0.025, 0.024, 0.022, 0.02, 0.019, 0.019, 0.02, 0.02, 0.021, 0.022, 0.024, 
    0.026, 0.028, 0.031, 0.034, 0.038, 0.043, 0.051, 0.057, 0.065, 0.073, 
    0.089, 0.114, 0.149, 0.202, 0.274, 0.357, 0.437, 0.498, 0.538, 0.564, 
    0.587, 0.622, 0.675, 0.741, 0.809, 0.874, 0.943, 1.02, 1.101, 1.173, 
    1.231, 1.271, 1.294, 1.291, 1.258, 1.202, 1.14, 1.093, 1.085, 1.122, 
    1.169, 1.195, 1.208, 1.233, 1.27, 1.3, 1.317, 1.315, 1.309, 1.309, 1.291, 
    1.207, 1.207 ;

 idx_rfr_Fe2O3_oray_roush_rl_ee = 0.158, 0.169, 0.184, 0.201, 0.23, 0.251, 
    0.224, 0.266, 0.348, 0.452, 0.737, 0.857, 0.938, 0.648, 0.381, 0.25, 
    0.18, 0.134, 0.114, 0.082, 0.05, 0.062, 0.092, 0.136, 0.221, 0.376, 
    0.479, 0.392, 0.249, 0.184, 0.145, 0.129, 0.121, 0.129, 0.2, 0.231, 
    0.189, 0.14, 0.103, 0.08, 0.067, 0.058, 0.051, 0.047, 0.044, 0.042, 
    0.041, 0.04, 0.039, 0.035, 0.029, 0.021, 0.016, 0.012, 0.01, 0.009, 
    0.009, 0.009, 0.009, 0.01, 0.011, 0.011, 0.012, 0.012, 0.013, 0.014, 
    0.014, 0.015, 0.015, 0.016, 0.016, 0.017, 0.017, 0.017, 0.018, 0.018, 
    0.018, 0.018, 0.019, 0.019, 0.019, 0.02, 0.02, 0.02, 0.021, 0.021, 0.021, 
    0.021, 0.021, 0.022, 0.022, 0.022, 0.022, 0.022, 0.023, 0.023, 0.023, 
    0.023, 0.023, 0.023, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.026, 
    0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.027, 
    0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 
    0.027, 0.027, 0.027, 0.027, 0.027, 0.028, 0.028, 0.028, 0.028, 0.028, 
    0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 
    0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.029, 0.029, 0.029, 
    0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 
    0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 
    0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 
    0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 
    0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 
    0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 
    0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.033, 0.033, 
    0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 
    0.033, 0.033, 0.033, 0.033, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 
    0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.035, 0.035, 0.035, 0.035, 
    0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.036, 0.036, 0.036, 0.036, 
    0.036, 0.036, 0.037, 0.037, 0.037, 0.038, 0.038, 0.038, 0.039, 0.039, 
    0.039, 0.04, 0.04, 0.041, 0.042, 0.042, 0.043, 0.044, 0.045, 0.047, 
    0.048, 0.05, 0.052, 0.054, 0.056, 0.058, 0.058, 0.058, 0.059, 0.059, 
    0.061, 0.063, 0.065, 0.068, 0.07, 0.072, 0.075, 0.078, 0.08, 0.082, 
    0.083, 0.082, 0.081, 0.078, 0.074, 0.07, 0.067, 0.067, 0.069, 0.072, 
    0.073, 0.073, 0.074, 0.076, 0.077, 0.077, 0.077, 0.076, 0.075, 0.077, 
    0.075, 0.075 ;

 idx_rfr_Fe2O3_oray_roush_img_ee = 0.016, 0.017, 0.013, 0.009, 0.004, 0.083, 
    0.072, 0.017, 0.053, 0.116, 0.368, 1.237, 1.033, 0.655, 0.443, 0.328, 
    0.256, 0.191, 0.12, 0.032, 0.051, 0.053, 0.066, 0.098, 0.174, 0.423, 
    0.481, 0.41, 0.305, 0.242, 0.195, 0.137, 0.069, 0.071, 0.138, 0.211, 
    0.22, 0.203, 0.18, 0.16, 0.143, 0.13, 0.118, 0.107, 0.096, 0.087, 0.077, 
    0.065, 0.051, 0.034, 0.016, 0.004, 0.009, 0.011, 0.011, 0.01, 0.01, 
    0.009, 0.008, 0.008, 0.007, 0.007, 0.007, 0.007, 0.006, 0.006, 0.006, 
    0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.005, 0.005, 
    0.005, 0.005, 0.005, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.003, 0.003, 0.002, 0.002, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.002, 0.002, 0.002, 0.002, 
    0.003, 0.003, 0.003, 0.002, 0.002, 0.002, 0.003, 0.003, 0.002, 0.002, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.002, 0.003, 
    0.002, 0.002, 0.002, 0.003, 0.003, 0.003, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.003, 0.003, 0.002, 0.002, 0.002, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.003, 0.003, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.002, 0.002, 0.002, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.003, 0.003, 0.003, 0.004, 0.004, 
    0.005, 0.005, 0.006, 0.008, 0.01, 0.013, 0.017, 0.024, 0.031, 0.037, 
    0.042, 0.045, 0.047, 0.048, 0.051, 0.055, 0.06, 0.064, 0.068, 0.072, 
    0.076, 0.079, 0.08, 0.08, 0.079, 0.076, 0.072, 0.068, 0.064, 0.062, 
    0.061, 0.061, 0.062, 0.062, 0.06, 0.058, 0.057, 0.054, 0.05, 0.044, 
    0.038, 0.031, 0.023, 0.029, 0.039, 0.039 ;

 idx_rfr_Fe2O3_oray_roush_nr = 0.49191, 0.50341, 0.51795, 0.5325, 0.5545, 
    0.5686, 0.5503, 0.57785, 0.61915, 0.65705, 0.7238, 0.8026, 0.85685, 
    0.8886, 0.8962, 0.87885, 0.8455, 0.76735, 0.55465, 0.2673, 0.2136, 
    0.30055, 0.38405, 0.4589, 0.54725, 0.66285, 0.7658, 0.8232, 0.83235, 
    0.8041, 0.7558, 0.5983, 0.40755, 0.432, 0.56715, 0.6719, 0.742, 0.7914, 
    0.82, 0.827, 0.81525, 0.7938, 0.76545, 0.71965, 0.6524, 0.5648, 0.4592, 
    0.3196, 0.17695, 0.0797, 0.03555, 0.0216, 0.0189, 0.02125, 0.0264, 
    0.03295, 0.04045, 0.04805, 0.0557, 0.06315, 0.06995, 0.07605, 0.0818, 
    0.08715, 0.0921, 0.09705, 0.10145, 0.10555, 0.10935, 0.11295, 0.1166, 
    0.1199, 0.1228, 0.12515, 0.1272, 0.1294, 0.1317, 0.1339, 0.136, 0.1381, 
    0.1403, 0.14235, 0.14425, 0.1461, 0.14785, 0.1493, 0.1507, 0.15205, 
    0.15345, 0.15485, 0.1562, 0.1575, 0.15885, 0.1601, 0.16125, 0.1624, 
    0.16345, 0.16425, 0.16525, 0.16615, 0.16705, 0.1679, 0.16875, 0.16955, 
    0.17035, 0.1712, 0.172, 0.17275, 0.17345, 0.1741, 0.1748, 0.17545, 
    0.17615, 0.1769, 0.17755, 0.1782, 0.17885, 0.1795, 0.1802, 0.1808, 
    0.1813, 0.1819, 0.18245, 0.18295, 0.1835, 0.18395, 0.1844, 0.18485, 
    0.1853, 0.1857, 0.186, 0.18635, 0.1868, 0.18725, 0.1876, 0.18785, 0.1881, 
    0.18845, 0.18875, 0.189, 0.1892, 0.18945, 0.18975, 0.1901, 0.19045, 
    0.19075, 0.1911, 0.19135, 0.1915, 0.1917, 0.19195, 0.19225, 0.1925, 
    0.19275, 0.19295, 0.1932, 0.19345, 0.19365, 0.19385, 0.194, 0.19415, 
    0.19435, 0.19455, 0.19475, 0.19495, 0.1951, 0.1953, 0.19545, 0.19565, 
    0.19585, 0.19605, 0.19615, 0.1963, 0.19645, 0.19665, 0.19685, 0.19695, 
    0.1971, 0.1972, 0.1974, 0.1975, 0.19765, 0.19775, 0.1979, 0.19795, 
    0.19815, 0.19825, 0.1984, 0.19855, 0.19865, 0.1988, 0.19885, 0.199, 
    0.1991, 0.19925, 0.1993, 0.1994, 0.19955, 0.1997, 0.1998, 0.19985, 
    0.19995, 0.20005, 0.20015, 0.20025, 0.2003, 0.2004, 0.2005, 0.20055, 
    0.20065, 0.20075, 0.20085, 0.20095, 0.2011, 0.20125, 0.2014, 0.20155, 
    0.20165, 0.20175, 0.20175, 0.20165, 0.2016, 0.2018, 0.20205, 0.2022, 
    0.2022, 0.20225, 0.20235, 0.20245, 0.20255, 0.20265, 0.2027, 0.2028, 
    0.2028, 0.2029, 0.20295, 0.20305, 0.20305, 0.20315, 0.2032, 0.20325, 
    0.2033, 0.20335, 0.2034, 0.20345, 0.20355, 0.2036, 0.2037, 0.20375, 
    0.2038, 0.20385, 0.2039, 0.20395, 0.20405, 0.2041, 0.20415, 0.2042, 
    0.20425, 0.20435, 0.20435, 0.20435, 0.20435, 0.2044, 0.2045, 0.2046, 
    0.20465, 0.2047, 0.20475, 0.2048, 0.2049, 0.20495, 0.20495, 0.205, 
    0.20505, 0.2051, 0.20515, 0.2051, 0.20515, 0.20515, 0.20515, 0.20515, 
    0.2052, 0.2052, 0.2051, 0.2051, 0.20525, 0.2053, 0.2053, 0.20535, 
    0.20545, 0.2055, 0.2055, 0.2055, 0.2055, 0.20555, 0.20555, 0.2056, 
    0.20565, 0.2057, 0.20575, 0.2058, 0.20585, 0.20585, 0.2059, 0.206, 
    0.20605, 0.2061, 0.20615, 0.2062, 0.2062, 0.20615, 0.20615, 0.20625, 
    0.2063, 0.20635, 0.20635, 0.20635, 0.2064, 0.20645, 0.2064, 0.20635, 
    0.20635, 0.2064, 0.20645, 0.20645, 0.20655, 0.20655, 0.2066, 0.20665, 
    0.20665, 0.20665, 0.2067, 0.20675, 0.20675, 0.20675, 0.20685, 0.2069, 
    0.20695, 0.207, 0.20705, 0.20705, 0.2071, 0.20715, 0.2072, 0.2072, 
    0.20715, 0.20715, 0.2072, 0.20725, 0.2073, 0.2073, 0.20735, 0.20735, 
    0.20735, 0.2074, 0.2075, 0.2076, 0.2076, 0.2075, 0.2074, 0.2074, 0.2075, 
    0.2076, 0.2076, 0.2076, 0.2077, 0.2077, 0.20765, 0.2076, 0.2076, 0.2076, 
    0.2076, 0.20755, 0.2075, 0.2075, 0.2075, 0.20745, 0.2074, 0.2074, 0.2074, 
    0.20745, 0.2075, 0.2075, 0.20755, 0.20765, 0.2077, 0.20775, 0.20775, 
    0.2077, 0.2077, 0.2077, 0.20775, 0.20775, 0.20775, 0.20775, 0.20775, 
    0.20785, 0.2079, 0.2079, 0.2079, 0.2079, 0.20795, 0.208, 0.208, 0.208, 
    0.208, 0.20805, 0.20805, 0.20805, 0.20805, 0.2081, 0.2081, 0.2081, 
    0.2081, 0.20815, 0.20815, 0.20815, 0.20815, 0.2082, 0.2082, 0.2082, 
    0.20825, 0.20825, 0.2083, 0.20835, 0.20835, 0.20835, 0.20835, 0.2084, 
    0.2084, 0.2084, 0.2084, 0.20845, 0.2085, 0.20855, 0.2086, 0.20865, 
    0.2087, 0.2087, 0.2087, 0.2087, 0.2087, 0.2087, 0.2086, 0.2084, 0.2083, 
    0.20825, 0.2084, 0.20855, 0.20865, 0.2088, 0.20895, 0.20915, 0.2093, 
    0.20935, 0.2093, 0.20935, 0.2094, 0.20945, 0.2095, 0.20955, 0.2096, 
    0.2097, 0.2098, 0.20985, 0.2099, 0.20995, 0.21, 0.21, 0.21005, 0.2101, 
    0.2101, 0.21015, 0.21025, 0.2104, 0.21055, 0.2107, 0.21075, 0.21075, 
    0.2108, 0.2109, 0.211, 0.2111, 0.2112, 0.2113, 0.21145, 0.2116, 0.21175, 
    0.2119, 0.212, 0.21205, 0.21215, 0.21225, 0.2124, 0.21255, 0.21275, 
    0.21295, 0.21315, 0.21335, 0.21355, 0.21365, 0.2138, 0.21395, 0.21415, 
    0.2144, 0.2147, 0.21495, 0.2152, 0.21535, 0.21555, 0.21575, 0.216, 
    0.21625, 0.21645, 0.2167, 0.217, 0.2174, 0.21775, 0.21805, 0.2183, 
    0.2185, 0.2188, 0.2191, 0.21945, 0.21985, 0.2202, 0.22055, 0.221, 
    0.22145, 0.22185, 0.22225, 0.22265, 0.2231, 0.2236, 0.224, 0.2244, 
    0.2247, 0.225, 0.22535, 0.2257, 0.22615, 0.22665, 0.2272, 0.22765, 
    0.22815, 0.2286, 0.2291, 0.22965, 0.2302, 0.23085, 0.2315, 0.23235, 
    0.2334, 0.2346, 0.23585, 0.2371, 0.23845, 0.2399, 0.2415, 0.24315, 
    0.2449, 0.2467, 0.2487, 0.2509, 0.25325, 0.2559, 0.25865, 0.2615, 0.2649, 
    0.269, 0.2739, 0.27925, 0.2852, 0.2913, 0.29665, 0.3001, 0.30095, 0.2998, 
    0.2979, 0.2967, 0.29735, 0.3, 0.30365, 0.3069, 0.30915, 0.311, 0.31315, 
    0.31535, 0.31665, 0.3162, 0.31395, 0.3099, 0.30375, 0.29475, 0.2828, 
    0.26965, 0.25845, 0.25225, 0.253, 0.258, 0.2609, 0.25975, 0.25775, 
    0.2582, 0.2596, 0.2595, 0.2573, 0.2527, 0.2484, 0.24695, 0.2455, 0.23995, 
    0.23995 ;

}

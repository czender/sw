// ncgen -b -o ~ammann/DATA/AERO/idx_rfr/idx_rfr_NNM98.nc ~ammann/DATA/AERO/idx_rfr/idx_rfr_NNM98.cdl
// ncks -C -H -s %9.5f -v bnd,idx_rfr_H2SO4_210K_61_NNM98_img,idx_rfr_H2SO4_210K_61_NNM98_rl,idx_rfr_H2SO4_220K_72_NNM98_img,idx_rfr_H2SO4_220K_72_NNM98_rl /ammann/DATA/AERO/idx_rfr/idx_rfr_NNM98.nc

netcdf idx_rfr_NNM98 {
dimensions:
        bnd=2112;
        bnd_PaW75=227;
        bnd_HSL88=57;
variables:
        :history = "";
        :source="
Caspar Ammann : Thu Jun 18 MDT 1999:
HSL88 : from /home/zender/idx_rfr/hitran/shettle.dat
HSL88 : Hummel, J. R., Shettle, E. P. and Longtin, D. R. (1988) 
        A New Background Stratospheric Aerosol Model for Use in 
        Atmospheric Radiation Models, AFGL-TR-88-0166, 
        Air Force Geophysics Laboratory, Hanscom AFB, MA, August 1988.
HSL88 : Range used : 0.2 - 0.337 micron
HSL88 : optical constants for H2SO4 75% for 215.
NNM98 = Niedziela, Norman, Miller and Worsnop, 1998: Temperature- and 
        composition-dependent infrared optical constants for sulfuric 
        acid. GRL 25, 4477-4480.  
        Optical constants calculated for different temperatures and 
        mixing ratios H2SO4 with Water Copied from frenchie.chem.unc.edu
Range:  2.12--12.11 micron, these indices are also shown graphically in NNM98.
PaW75 : Kent F. Palmer and Dudley Williams, 1975: Optical constants of 
        sulfuric acid; application to the clouds of Venus? 
        Applied Optics 14, 1, p. 208-219.  
        Calculated for 300K and different mixing ratios H2SO4 with Water. 
        Selected 75% H2SO4 25%. Copied from palmer_w.dat in 
        /home/zender/idx_rfr/hitran
Range:  0.36--25.0 microns, these indices are also shown graphically in PaW75.

Caspar Ammann : Thu Apr 6 2001: Fix of NNM98 data below 2.1 micron.";

        float bnd(bnd);
        bnd:long_name = "Band center wavelength";
        bnd:units = "micron";
        bnd:C_format = "%.7g";

        float bnd_PaW75(bnd_PaW75);
        bnd_PaW75:long_name = "Band center wavelength";
        bnd_PaW75:units = "micron";
        bnd_PaW75:C_format = "%.3g";

        float bnd_HSL88(bnd_HSL88);
        bnd_HSL88:long_name = "Band center wavelength";
        bnd_HSL88:units = "micron";
        bnd_HSL88:C_format = "%.3g";

        float idx_rfr_H2SO4_210K_61_NNM98_rl(bnd);
        idx_rfr_H2SO4_210K_61_NNM98_rl:long_name = "Sulfate 61% real index of refraction";
        idx_rfr_H2SO4_210K_61_NNM98_rl:units = "";
        idx_rfr_H2SO4_210K_61_NNM98_rl:C_format = "%.5g";

        float idx_rfr_H2SO4_210K_61_NNM98_img(bnd);
        idx_rfr_H2SO4_210K_61_NNM98_img:long_name = "Sulfate 61% imaginary index of refraction";
        idx_rfr_H2SO4_210K_61_NNM98_img:units = "";
        idx_rfr_H2SO4_210K_61_NNM98_img:C_format = "%.6g";

        float idx_rfr_H2SO4_220K_72_NNM98_rl(bnd);
        idx_rfr_H2SO4_220K_72_NNM98_rl:long_name = "Sulfate 72% real index of refraction";
        idx_rfr_H2SO4_220K_72_NNM98_rl:units = "";
        idx_rfr_H2SO4_220K_72_NNM98_rl:C_format = "%.5g";

        float idx_rfr_H2SO4_220K_72_NNM98_img(bnd);
        idx_rfr_H2SO4_220K_72_NNM98_img:long_name = "Sulfate 72% imaginary index of refraction";
        idx_rfr_H2SO4_220K_72_NNM98_img:units = "";
        idx_rfr_H2SO4_220K_72_NNM98_img:C_format = "%.6g";

        float idx_rfr_H2SO4_300K_PaW75_rl(bnd_PaW75);
        idx_rfr_H2SO4_300K_PaW75_rl:long_name = "Sulfate 75% real index of refraction";
        idx_rfr_H2SO4_300K_PaW75_rl:units = "";
        idx_rfr_H2SO4_300K_PaW75_rl:C_format = "%.3g";

        float idx_rfr_H2SO4_300K_PaW75_img(bnd_PaW75);
        idx_rfr_H2SO4_300K_PaW75_img:long_name = "Sulfate 75% imaginary index of refraction";
        idx_rfr_H2SO4_300K_PaW75_img:units = "";
        idx_rfr_H2SO4_300K_PaW75_img:C_format = "%.6g";

        float idx_rfr_H2SO4_215K_75_HSL88_rl(bnd_HSL88);
        idx_rfr_H2SO4_215K_75_HSL88_rl:long_name = "Sulfate 75% real index of refraction";
        idx_rfr_H2SO4_215K_75_HSL88_rl:units = "";
        idx_rfr_H2SO4_215K_75_HSL88_rl:C_format = "%.3g";

        float idx_rfr_H2SO4_215K_75_HSL88_img(bnd_HSL88);
        idx_rfr_H2SO4_215K_75_HSL88_img:long_name = "Sulfate 75% imaginary index of refraction";
        idx_rfr_H2SO4_215K_75_HSL88_img:units = "";
        idx_rfr_H2SO4_215K_75_HSL88_img:C_format = "%.5g";


data:

 bnd = 
0.2, 0.25, 0.3, 0.337,
0.360,  0.445,  0.449,  0.556,  0.702,  0.714,  0.725,  0.735,  0.746,  0.758,
0.769,  0.781,  0.794,  0.806,  0.820,  0.833,  0.847,  0.862,  0.877,  0.893,  
0.909,  0.926,  0.943,  0.962,  0.980,  1.000,  1.020,  1.042,  1.064,  1.087,  
1.111,  1.136,  1.163,  1.190,  1.220,  1.250,  1.266,  1.282,  1.299,  1.316,  
1.333,  1.351,  1.370,  1.389,  1.408,  1.429,  1.449,  1.471,  1.493,  1.515,  
1.538,  1.562,  1.587,  1.613,  1.639,  1.667,  1.695,  1.724,  1.754,  1.786,  
1.818,  1.852,  1.887,  1.923,  1.961,  2.000,  2.041,  2.083,
2.1272879,  2.1281612,  2.1290352,  2.1299098,  2.1307852,  2.1316614,  2.1325383,  2.1334159,  2.1342943,  2.1351731,  2.1360531,  2.1369333,  2.1378148,  2.1386967,  2.1395793,  2.1404626,  2.1413469,  2.1422317,  2.1431172,  2.1440036,  2.1448905,  2.1457784,  2.1466668,  2.1475563,  2.1484461,  2.1493371,  2.1502283,  2.1511207,  2.1520135,  2.1529074,  2.1538017,  2.1546967,  2.1555929,  2.1564894,  2.1573870,  2.1582849,  2.1591840,  2.1600835,  2.1609840,  2.1618850,  2.1627872,  2.1636896,  2.1645932,  2.1654973,  2.1664023,  2.1673081,  2.1682143,  2.1691215,  2.1700294,  2.1709383,  2.1718476,  2.1727579,  2.1736689,  2.1745808,  2.1754932,  2.1764066,  2.1773207,  2.1782355,  2.1791511,  2.1800673,  2.1809847,  2.1819024,  2.1828213,  2.1837406,  2.1846609,  2.1855819,  2.1865039,  2.1874263,  2.1883497,  2.1892738,  2.1901989,  2.1911244,  2.1920509,  2.1929784,  2.1939061,  2.1948352,  2.1957648,  2.1966951,  2.1976264,  2.1985583,  2.1994910,  2.2004247,  2.2013590,  2.2022943,  2.2032301,  2.2041669,  2.2051044,  2.2060428,  2.2069819,  2.2079217,  2.2088625,  2.2098041,  2.2107465,  2.2116895,  2.2126336,  2.2135782,  2.2145240,  2.2154703,  2.2164176,  2.2173655,  2.2183144,  2.2192640,  2.2202141,  2.2211657,  2.2221177,  2.2230706,  2.2240243,  2.2249789,  2.2259340,  2.2268903,  2.2278471,  2.2288051,  2.2297637,  2.2307231,  2.2316833,  2.2326446,  2.2336066,  2.2345691,  2.2355330,  2.2364972,  2.2374625,  2.2384284,  2.2393956,  2.2403634,  2.2413321,  2.2423012,  2.2432716,  2.2442427,  2.2452147,  2.2461874,  2.2471609,  2.2481356,  2.2491107,  2.2500870,  2.2510641,  2.2520421,  2.2530208,  2.2540002,  2.2549806,  2.2559621,  2.2569439,  2.2579272,  2.2589109,  2.2598958,  2.2608812,  2.2618675,  2.2628551,  2.2638428,  2.2648323,  2.2658219,  2.2668126,  2.2678041,  2.2687969,  2.2697899,  2.2707844,  2.2717793,  2.2727754,  2.2737720,  2.2747698,  2.2757685,  2.2767677,  2.2777681,  2.2787695,  2.2797716,  2.2807746,  2.2817783,  2.2827830,  2.2837889,  2.2847953,  2.2858028,  2.2868109,  2.2878203,  2.2888303,  2.2898412,  2.2908533,  2.2918656,  2.2928796,  2.2938938,  2.2949095,  2.2959259,  2.2969432,  2.2979612,  2.2989805,  2.3000002,  2.3010211,  2.3020430,  2.3030653,  2.3040891,  2.3051136,  2.3061390,  2.3071654,  2.3081927,  2.3092208,  2.3102498,  2.3112798,  2.3123109,  2.3133423,  2.3143754,  2.3154089,  2.3164437,  2.3174789,  2.3185153,  2.3195529,  2.3205910,  2.3216302,  2.3226705,  2.3237116,  2.3247535,  2.3257966,  2.3268404,  2.3278854,  2.3289311,  2.3299778,  2.3310254,  2.3320739,  2.3331234,  2.3341739,  2.3352253,  2.3362777,  2.3373313,  2.3383853,  2.3394406,  2.3404968,  2.3415542,  2.3426120,  2.3436713,  2.3447311,  2.3457921,  2.3468540,  2.3479168,  2.3489807,  2.3500454,  2.3511114,  2.3521781,  2.3532460,  2.3543146,  2.3553841,  2.3564548,  2.3575265,  2.3585989,  2.3596725,  2.3607471,  2.3618224,  2.3628991,  2.3639765,  2.3650551,  2.3661342,  2.3672149,  2.3682961,  2.3693788,  2.3704619,  2.3715465,  2.3726318,  2.3737183,  2.3748055,  2.3758941,  2.3769834,  2.3780735,  2.3791652,  2.3802571,  2.3813508,  2.3824449,  2.3835406,  2.3846366,  2.3857343,  2.3868327,  2.3879323,  2.3890324,  2.3901341,  2.3912363,  2.3923397,  2.3934445,  2.3945498,  2.3956566,  2.3967638,  2.3978727,  2.3989823,  2.4000928,  2.4012043,  2.4023173,  2.4034309,  2.4045458,  2.4056616,  2.4067786,  2.4078963,  2.4090149,  2.4101350,  2.4112561,  2.4123781,  2.4135010,  2.4146254,  2.4157503,  2.4168768,  2.4180038,  2.4191325,  2.4202616,  2.4213922,  2.4225235,  2.4236562,  2.4247897,  2.4259243,  2.4270601,  2.4281969,  2.4293349,  2.4304738,  2.4316139,  2.4327548,  2.4338970,  2.4350400,  2.4361846,  2.4373298,  2.4384763,  2.4396238,  2.4407723,  2.4419219,  2.4430728,  2.4442246,  2.4453778,  2.4465318,  2.4476869,  2.4488428,  2.4500003,  2.4511588,  2.4523182,  2.4534788,  2.4546404,  2.4558032,  2.4569671,  2.4581323,  2.4592981,  2.4604654,  2.4616337,  2.4628031,  2.4639738,  2.4651451,  2.4663179,  2.4674921,  2.4686670,  2.4698429,  2.4710202,  2.4721987,  2.4733782,  2.4745588,  2.4757407,  2.4769235,  2.4781075,  2.4792924,  2.4804788,  2.4816661,  2.4828544,  2.4840443,  2.4852352,  2.4864271,  2.4876201,  2.4888144,  2.4900100,  2.4912064,  2.4924040,  2.4936030,  2.4948030,  2.4960041,  2.4972064,  2.4984100,  2.4996145,  2.5008202,  2.5020273,  2.5032353,  2.5044446,  2.5056553,  2.5068669,  2.5080795,  2.5092936,  2.5105085,  2.5117252,  2.5129426,  2.5141613,  2.5153811,  2.5166020,  2.5178244,  2.5190477,  2.5202725,  2.5214982,  2.5227253,  2.5239534,  2.5251827,  2.5264137,  2.5276453,  2.5288785,  2.5301127,  2.5313478,  2.5325844,  2.5338223,  2.5350611,  2.5363016,  2.5375433,  2.5387857,  2.5400295,  2.5412748,  2.5425210,  2.5437689,  2.5450172,  2.5462677,  2.5475187,  2.5487711,  2.5500247,  2.5512795,  2.5525360,  2.5537932,  2.5550520,  2.5563118,  2.5575731,  2.5588355,  2.5600989,  2.5613637,  2.5626302,  2.5638976,  2.5651662,  2.5664361,  2.5677071,  2.5689795,  2.5702529,  2.5715280,  2.5728042,  2.5740817,  2.5753603,  2.5766404,  2.5779219,  2.5792041,  2.5804882,  2.5817730,  2.5830595,  2.5843475,  2.5856361,  2.5869262,  2.5882180,  2.5895107,  2.5908051,  2.5921004,  2.5933969,  2.5946949,  2.5959942,  2.5972948,  2.5985968,  2.5999000,  2.6012046,  2.6025105,  2.6038172,  2.6051257,  2.6064358,  2.6077466,  2.6090591,  2.6103730,  2.6116879,  2.6130042,  2.6143219,  2.6156409,  2.6169615,  2.6182830,  2.6196060,  2.6209307,  2.6222560,  2.6235831,  2.6249118,  2.6262414,  2.6275723,  2.6289048,  2.6302385,  2.6315739,  2.6329103,  2.6342483,  2.6355877,  2.6369281,  2.6382701,  2.6396136,  2.6409578,  2.6423039,  2.6436515,  2.6450005,  2.6463504,  2.6477020,  2.6490548,  2.6504092,  2.6517649,  2.6531219,  2.6544807,  2.6558404,  2.6572018,  2.6585646,  2.6599286,  2.6612937,  2.6626608,  2.6640291,  2.6653986,  2.6667697,  2.6681423,  2.6695163,  2.6708918,  2.6722684,  2.6736465,  2.6750262,  2.6764071,  2.6777897,  2.6791735,  2.6805584,  2.6819453,  2.6833336,  2.6847234,  2.6861141,  2.6875067,  2.6889005,  2.6902962,  2.6916928,  2.6930912,  2.6944909,  2.6958921,  2.6972947,  2.6986990,  2.7001045,  2.7015116,  2.7029200,  2.7043300,  2.7057414,  2.7071543,  2.7085686,  2.7099845,  2.7114019,  2.7128208,  2.7142413,  2.7156630,  2.7170861,  2.7185111,  2.7199371,  2.7213650,  2.7227943,  2.7242250,  2.7256575,  2.7270913,  2.7285266,  2.7299635,  2.7314017,  2.7328415,  2.7342830,  2.7357261,  2.7371705,  2.7386162,  2.7400637,  2.7415128,  2.7429633,  2.7444153,  2.7458689,  2.7473242,  2.7487807,  2.7502389,  2.7516987,  2.7531600,  2.7546232,  2.7560875,  2.7575536,  2.7590210,  2.7604902,  2.7619607,  2.7634332,  2.7649069,  2.7663822,  2.7678592,  2.7693381,  2.7708180,  2.7722995,  2.7737830,  2.7752678,  2.7767546,  2.7782426,  2.7797322,  2.7812235,  2.7827163,  2.7842107,  2.7857070,  2.7872045,  2.7887039,  2.7902050,  2.7917073,  2.7932117,  2.7947176,  2.7962248,  2.7977338,  2.7992446,  2.8007567,  2.8022704,  2.8037858,  2.8053033,  2.8068221,  2.8083427,  2.8098648,  2.8113887,  2.8129141,  2.8144412,  2.8159699,  2.8175001,  2.8190324,  2.8205662,  2.8221016,  2.8236384,  2.8251772,  2.8267176,  2.8282599,  2.8298039,  2.8313494,  2.8328965,  2.8344452,  2.8359959,  2.8375480,  2.8391023,  2.8406579,  2.8422153,  2.8437743,  2.8453350,  2.8468974,  2.8484616,  2.8500278,  2.8515954,  2.8531649,  2.8547359,  2.8563087,  2.8578835,  2.8594599,  2.8610377,  2.8626175,  2.8641994,  2.8657825,  2.8673675,  2.8689544,  2.8705428,  2.8721333,  2.8737254,  2.8753190,  2.8769147,  2.8785124,  2.8801115,  2.8817122,  2.8833151,  2.8849194,  2.8865261,  2.8881340,  2.8897438,  2.8913555,  2.8929691,  2.8945844,  2.8962014,  2.8978205,  2.8994408,  2.9010634,  2.9026880,  2.9043140,  2.9059422,  2.9075718,  2.9092035,  2.9108372,  2.9124720,  2.9141092,  2.9157484,  2.9173892,  2.9190319,  2.9206762,  2.9223225,  2.9239709,  2.9256213,  2.9272733,  2.9289269,  2.9305825,  2.9322402,  2.9338996,  2.9355607,  2.9372241,  2.9388890,  2.9405560,  2.9422250,  2.9438958,  2.9455683,  2.9472430,  2.9489195,  2.9505978,  2.9522784,  2.9539604,  2.9556448,  2.9573307,  2.9590187,  2.9607086,  2.9624004,  2.9640939,  2.9657898,  2.9674873,  2.9691870,  2.9708884,  2.9725921,  2.9742973,  2.9760048,  2.9777145,  2.9794257,  2.9811392,  2.9828541,  2.9845712,  2.9862905,  2.9880116,  2.9897349,  2.9914603,  2.9931872,  2.9949167,  2.9966476,  2.9983809,  3.0001159,  3.0018532,  3.0035925,  3.0053337,  3.0070770,  3.0088222,  3.0105691,  3.0123186,  3.0140700,  3.0158234,  3.0175788,  3.0193365,  3.0210958,  3.0228574,  3.0246210,  3.0263867,  3.0281546,  3.0299244,  3.0316963,  3.0334702,  3.0352461,  3.0370243,  3.0388045,  3.0405869,  3.0423713,  3.0441577,  3.0459464,  3.0477369,  3.0495296,  3.0513248,  3.0531216,  3.0549209,  3.0567222,  3.0585253,  3.0603309,  3.0621386,  3.0639482,  3.0657601,  3.0675743,  3.0693903,  3.0712087,  3.0730295,  3.0748520,  3.0766768,  3.0785038,  3.0803332,  3.0821645,  3.0839980,  3.0858335,  3.0876713,  3.0895116,  3.0913539,  3.0931985,  3.0950451,  3.0968940,  3.0987451,  3.1005983,  3.1024539,  3.1043117,  3.1061718,  3.1080341,  3.1098983,  3.1117649,  3.1136341,  3.1155050,  3.1173785,  3.1192544,  3.1211321,  3.1230125,  3.1248949,  3.1267796,  3.1286666,  3.1305559,  3.1324477,  3.1343415,  3.1362371,  3.1381359,  3.1400368,  3.1419396,  3.1438448,  3.1457527,  3.1476629,  3.1495750,  3.1514897,  3.1534066,  3.1553261,  3.1572475,  3.1591716,  3.1610980,  3.1630263,  3.1649575,  3.1668909,  3.1688268,  3.1707649,  3.1727052,  3.1746480,  3.1765935,  3.1785412,  3.1804910,  3.1824436,  3.1843984,  3.1863558,  3.1883154,  3.1902771,  3.1922417,  3.1942086,  3.1961777,  3.1981494,  3.2001235,  3.2021003,  3.2040794,  3.2060611,  3.2080448,  3.2100315,  3.2120202,  3.2140117,  3.2160053,  3.2180016,  3.2200003,  3.2220016,  3.2240052,  3.2260115,  3.2280202,  3.2300315,  3.2320452,  3.2340615,  3.2360802,  3.2381015,  3.2401254,  3.2421520,  3.2441807,  3.2462118,  3.2482460,  3.2502823,  3.2523212,  3.2543633,  3.2564073,  3.2584541,  3.2605035,  3.2625554,  3.2646098,  3.2666671,  3.2687268,  3.2707891,  3.2728541,  3.2749214,  3.2769914,  3.2790642,  3.2811394,  3.2832174,  3.2852981,  3.2873816,  3.2894673,  3.2915559,  3.2936471,  3.2957411,  3.2978377,  3.2999368,  3.3020384,  3.3041430,  3.3062501,  3.3083601,  3.3104727,  3.3125880,  3.3147063,  3.3168271,  3.3189504,  3.3210764,  3.3232055,  3.3253369,  3.3274715,  3.3296087,  3.3317485,  3.3338912,  3.3360362,  3.3381844,  3.3403354,  3.3424890,  3.3446453,  3.3468046,  3.3489666,  3.3511314,  3.3532991,  3.3554697,  3.3576429,  3.3598189,  3.3619978,  3.3641796,  3.3663638,  3.3685513,  3.3707416,  3.3729346,  3.3751304,  3.3773293,  3.3795309,  3.3817356,  3.3839428,  3.3861532,  3.3883662,  3.3905826,  3.3928015,  3.3950236,  3.3972480,  3.3994756,  3.4017065,  3.4039397,  3.4061763,  3.4084160,  3.4106581,  3.4129035,  3.4151521,  3.4174032,  3.4196572,  3.4219146,  3.4241748,  3.4264379,  3.4287040,  3.4309731,  3.4332452,  3.4355206,  3.4377985,  3.4400799,  3.4423642,  3.4446516,  3.4469419,  3.4492352,  3.4515319,  3.4538312,  3.4561336,  3.4584394,  3.4607477,  3.4630599,  3.4653745,  3.4676926,  3.4700136,  3.4723380,  3.4746652,  3.4769957,  3.4793291,  3.4816658,  3.4840059,  3.4863486,  3.4886951,  3.4910443,  3.4933965,  3.4957521,  3.4981110,  3.5004728,  3.5028381,  3.5052066,  3.5075781,  3.5099530,  3.5123308,  3.5147121,  3.5170965,  3.5194845,  3.5218754,  3.5242698,  3.5266669,  3.5290675,  3.5314715,  3.5338790,  3.5362895,  3.5387032,  3.5411208,  3.5435410,  3.5459647,  3.5483921,  3.5508225,  3.5532560,  3.5556931,  3.5581336,  3.5605772,  3.5630243,  3.5654747,  3.5679288,  3.5703859,  3.5728467,  3.5753107,  3.5777781,  3.5802491,  3.5827234,  3.5852010,  3.5876822,  3.5901668,  3.5926549,  3.5951459,  3.5976410,  3.6001391,  3.6026409,  3.6051464,  3.6076553,  3.6101675,  3.6126833,  3.6152027,  3.6177254,  3.6202519,  3.6227818,  3.6253152,  3.6278522,  3.6303923,  3.6329365,  3.6354840,  3.6380353,  3.6405902,  3.6431484,  3.6457105,  3.6482763,  3.6508455,  3.6534183,  3.6559949,  3.6585751,  3.6611586,  3.6637461,  3.6663368,  3.6689317,  3.6715300,  3.6741321,  3.6767378,  3.6793473,  3.6819606,  3.6845775,  3.6871979,  3.6898227,  3.6924508,  3.6950827,  3.6977179,  3.7003574,  3.7030003,  3.7056472,  3.7082977,  3.7109523,  3.7136106,  3.7162728,  3.7189386,  3.7216084,  3.7242820,  3.7269595,  3.7296407,  3.7323258,  3.7350152,  3.7377079,  3.7404041,  3.7431049,  3.7458093,  3.7485180,  3.7512305,  3.7539468,  3.7566671,  3.7593913,  3.7621195,  3.7648513,  3.7675877,  3.7703278,  3.7730718,  3.7758198,  3.7785716,  3.7813277,  3.7840879,  3.7868519,  3.7896202,  3.7923925,  3.7951686,  3.7979491,  3.8007336,  3.8035219,  3.8063147,  3.8091114,  3.8119123,  3.8147173,  3.8175263,  3.8203394,  3.8231566,  3.8259783,  3.8288038,  3.8316336,  3.8344679,  3.8373060,  3.8401484,  3.8429952,  3.8458462,  3.8487012,  3.8515608,  3.8544242,  3.8572922,  3.8601642,  3.8630404,  3.8659213,  3.8688061,  3.8716958,  3.8745892,  3.8774874,  3.8803895,  3.8832965,  3.8862073,  3.8891227,  3.8920424,  3.8949668,  3.8978953,  3.9008281,  3.9037654,  3.9067073,  3.9096534,  3.9126041,  3.9155593,  3.9185188,  3.9214830,  3.9244516,  3.9274249,  3.9304025,  3.9333844,  3.9363711,  3.9393623,  3.9423578,  3.9453580,  3.9483628,  3.9513724,  3.9543862,  3.9574051,  3.9604282,  3.9634559,  3.9664886,  3.9695258,  3.9725676,  3.9756141,  3.9786651,  3.9817209,  3.9847813,  3.9878464,  3.9909163,  3.9939911,  3.9970706,  4.0001545,  4.0032434,  4.0063372,  4.0094361,  4.0125394,  4.0156474,  4.0187602,  4.0218782,  4.0250006,  4.0281277,  4.0312600,  4.0343971,  4.0375390,  4.0406861,  4.0438380,  4.0469952,  4.0501566,  4.0533233,  4.0564952,  4.0596714,  4.0628533,  4.0660396,  4.0692315,  4.0724277,  4.0756292,  4.0788360,  4.0820475,  4.0852642,  4.0884862,  4.0917130,  4.0949450,  4.0981822,  4.1014242,  4.1046720,  4.1079245,  4.1111822,  4.1144452,  4.1177125,  4.1209860,  4.1242647,  4.1275482,  4.1308370,  4.1341310,  4.1374307,  4.1407351,  4.1440454,  4.1473603,  4.1506810,  4.1540070,  4.1573381,  4.1606750,  4.1640162,  4.1673636,  4.1707163,  4.1740742,  4.1774378,  4.1808066,  4.1841812,  4.1875610,  4.1909466,  4.1943369,  4.1977334,  4.2011352,  4.2045426,  4.2079554,  4.2113733,  4.2147970,  4.2182264,  4.2216616,  4.2251024,  4.2285485,  4.2320004,  4.2354579,  4.2389212,  4.2423902,  4.2458649,  4.2493448,  4.2528305,  4.2563224,  4.2598195,  4.2633228,  4.2668319,  4.2703462,  4.2738667,  4.2773933,  4.2809253,  4.2844634,  4.2880073,  4.2915568,  4.2951126,  4.2986741,  4.3022413,  4.3058147,  4.3093934,  4.3129787,  4.3165698,  4.3201671,  4.3237700,  4.3273792,  4.3309946,  4.3346162,  4.3382430,  4.3418765,  4.3455157,  4.3491616,  4.3528132,  4.3564711,  4.3601346,  4.3638048,  4.3674812,  4.3711638,  4.3748527,  4.3785477,  4.3822489,  4.3859568,  4.3896704,  4.3933902,  4.3971167,  4.4008493,  4.4045887,  4.4083338,  4.4120855,  4.4158435,  4.4196081,  4.4233789,  4.4271564,  4.4309406,  4.4347310,  4.4385281,  4.4423313,  4.4461412,  4.4499578,  4.4537807,  4.4576101,  4.4614463,  4.4652891,  4.4691381,  4.4729943,  4.4768567,  4.4807267,  4.4846025,  4.4884853,  4.4923749,  4.4962711,  4.5001740,  4.5040841,  4.5080004,  4.5119243,  4.5158544,  4.5197916,  4.5237350,  4.5276856,  4.5316439,  4.5356083,  4.5395799,  4.5435586,  4.5475440,  4.5515370,  4.5555363,  4.5595431,  4.5635567,  4.5675778,  4.5716057,  4.5756407,  4.5796824,  4.5837312,  4.5877876,  4.5918517,  4.5959225,  4.6000004,  4.6040859,  4.6081781,  4.6122780,  4.6163855,  4.6204996,  4.6246219,  4.6287508,  4.6328874,  4.6370306,  4.6411819,  4.6453409,  4.6495070,  4.6536808,  4.6578622,  4.6620507,  4.6662469,  4.6704507,  4.6746626,  4.6788812,  4.6831083,  4.6873426,  4.6915841,  4.6958337,  4.7000909,  4.7043562,  4.7086291,  4.7129097,  4.7171979,  4.7214942,  4.7257981,  4.7301102,  4.7344298,  4.7387576,  4.7430930,  4.7474365,  4.7517881,  4.7561469,  4.7605143,  4.7648897,  4.7692733,  4.7736654,  4.7780647,  4.7824726,  4.7868891,  4.7913132,  4.7957454,  4.8001857,  4.8046346,  4.8090916,  4.8135571,  4.8180299,  4.8225121,  4.8270020,  4.8315005,  4.8360076,  4.8405232,  4.8450470,  4.8495793,  4.8541203,  4.8586698,  4.8632278,  4.8677940,  4.8723693,  4.8769526,  4.8815446,  4.8861456,  4.8907557,  4.8953738,  4.9000006,  4.9046364,  4.9092808,  4.9139342,  4.9185963,  4.9232674,  4.9279475,  4.9326358,  4.9373341,  4.9420404,  4.9467564,  4.9514813,  4.9562149,  4.9609575,  4.9657087,  4.9704704,  4.9752402,  4.9800200,  4.9848080,  4.9896059,  4.9944129,  4.9992290,  5.0040545,  5.0088892,  5.0137339,  5.0185871,  5.0234504,  5.0283227,  5.0332041,  5.0380955,  5.0429964,  5.0479069,  5.0528274,  5.0577569,  5.0626955,  5.0676446,  5.0726032,  5.0775714,  5.0825496,  5.0875378,  5.0925355,  5.0975423,  5.1025591,  5.1075864,  5.1126237,  5.1176710,  5.1227274,  5.1277952,  5.1328721,  5.1379590,  5.1430559,  5.1481633,  5.1532807,  5.1584082,  5.1635461,  5.1686950,  5.1738524,  5.1790214,  5.1842008,  5.1893897,  5.1945896,  5.1998000,  5.2050209,  5.2102513,  5.2154932,  5.2207460,  5.2260084,  5.2312818,  5.2365661,  5.2418613,  5.2471662,  5.2524829,  5.2578096,  5.2631478,  5.2684965,  5.2738562,  5.2792273,  5.2846079,  5.2900009,  5.2954040,  5.3008184,  5.3062439,  5.3116808,  5.3171291,  5.3225875,  5.3280582,  5.3335395,  5.3390326,  5.3445368,  5.3500524,  5.3555794,  5.3611169,  5.3666673,  5.3722281,  5.3778009,  5.3833857,  5.3889818,  5.3945894,  5.4002090,  5.4058399,  5.4114828,  5.4171371,  5.4228039,  5.4284825,  5.4341722,  5.4398742,  5.4455886,  5.4513149,  5.4570532,  5.4628034,  5.4685659,  5.4743409,  5.4801273,  5.4859266,  5.4917378,  5.4975615,  5.5033975,  5.5092463,  5.5151072,  5.5209804,  5.5268664,  5.5327644,  5.5386763,  5.5445991,  5.5505357,  5.5564852,  5.5624471,  5.5684214,  5.5744090,  5.5804100,  5.5864234,  5.5924497,  5.5984893,  5.6045408,  5.6106067,  5.6166854,  5.6227775,  5.6288824,  5.6350002,  5.6411324,  5.6472769,  5.6534352,  5.6596079,  5.6657929,  5.6719918,  5.6782045,  5.6844306,  5.6906700,  5.6969233,  5.7031908,  5.7094717,  5.7157669,  5.7220755,  5.7283988,  5.7347350,  5.7410855,  5.7474508,  5.7538295,  5.7602229,  5.7666302,  5.7730522,  5.7794876,  5.7859383,  5.7924027,  5.7988815,  5.8053761,  5.8118844,  5.8184071,  5.8249440,  5.8314967,  5.8380637,  5.8446450,  5.8512425,  5.8578539,  5.8644805,  5.8711214,  5.8777781,  5.8844500,  5.8911366,  5.8978391,  5.9045568,  5.9112897,  5.9180374,  5.9248009,  5.9315796,  5.9383740,  5.9451842,  5.9520097,  5.9588513,  5.9657083,  5.9725809,  5.9794698,  5.9863744,  5.9932952,  6.0002317,  6.0071850,  6.0141540,  6.0211382,  6.0281401,  6.0351577,  6.0421915,  6.0492420,  6.0563092,  6.0633926,  6.0704923,  6.0776091,  6.0847425,  6.0918927,  6.0990591,  6.1062431,  6.1134443,  6.1206617,  6.1278963,  6.1351485,  6.1424174,  6.1497040,  6.1570077,  6.1643291,  6.1716671,  6.1790233,  6.1863971,  6.1937881,  6.2011967,  6.2086234,  6.2160683,  6.2235298,  6.2310100,  6.2385087,  6.2460251,  6.2535591,  6.2611117,  6.2686830,  6.2762718,  6.2838793,  6.2915053,  6.2991500,  6.3068132,  6.3144951,  6.3221960,  6.3299150,  6.3376536,  6.3454103,  6.3531871,  6.3609819,  6.3687968,  6.3766308,  6.3844833,  6.3923554,  6.4002471,  6.4081588,  6.4160895,  6.4240403,  6.4320107,  6.4400005,  6.4480104,  6.4560404,  6.4640903,  6.4721603,  6.4802508,  6.4883614,  6.4964919,  6.5046425,  6.5128145,  6.5210071,  6.5292196,  6.5374537,  6.5457082,  6.5539827,  6.5622787,  6.5705962,  6.5789347,  6.5872941,  6.5956755,  6.6040769,  6.6125002,  6.6209455,  6.6294127,  6.6379008,  6.6464109,  6.6549430,  6.6634970,  6.6720724,  6.6806707,  6.6892905,  6.6979332,  6.7065983,  6.7152858,  6.7239957,  6.7327275,  6.7414832,  6.7502608,  6.7590618,  6.7678857,  6.7767324,  6.7856030,  6.7944961,  6.8034129,  6.8123527,  6.8213162,  6.8303041,  6.8393145,  6.8483496,  6.8574080,  6.8664904,  6.8755970,  6.8847284,  6.8938837,  6.9030638,  6.9122672,  6.9214954,  6.9307489,  6.9400272,  6.9493303,  6.9586582,  6.9680119,  6.9773903,  6.9867930,  6.9962220,  7.0056763,  7.0151563,  7.0246615,  7.0341930,  7.0437508,  7.0533338,  7.0629430,  7.0725789,  7.0822415,  7.0919294,  7.1016450,  7.1113863,  7.1211543,  7.1309495,  7.1407719,  7.1506214,  7.1604981,  7.1704021,  7.1803336,  7.1902919,  7.2002783,  7.2102928,  7.2203350,  7.2304053,  7.2405038,  7.2506304,  7.2607846,  7.2709680,  7.2811804,  7.2914209,  7.3016911,  7.3119898,  7.3223171,  7.3326735,  7.3430600,  7.3534756,  7.3639212,  7.3743958,  7.3849015,  7.3954358,  7.4060006,  7.4165955,  7.4272213,  7.4378772,  7.4485641,  7.4592814,  7.4700303,  7.4808083,  7.4916186,  7.5024610,  7.5133343,  7.5242391,  7.5351753,  7.5461435,  7.5571432,  7.5681758,  7.5792403,  7.5903373,  7.6014671,  7.6126294,  7.6238246,  7.6350527,  7.6463132,  7.6576076,  7.6689358,  7.6802969,  7.6916924,  7.7031217,  7.7145844,  7.7260809,  7.7376122,  7.7491784,  7.7607789,  7.7724147,  7.7840848,  7.7957907,  7.8075309,  7.8193069,  7.8311186,  7.8429661,  7.8548498,  7.8667688,  7.8787246,  7.8907161,  7.9027448,  7.9148102,  7.9269118,  7.9390516,  7.9512281,  7.9634418,  7.9756927,  7.9879823,  8.0003090,  8.0126743,  8.0250788,  8.0375204,  8.0500011,  8.0625200,  8.0750780,  8.0876760,  8.1003132,  8.1129904,  8.1257067,  8.1384630,  8.1512585,  8.1640949,  8.1769724,  8.1898899,  8.2028484,  8.2158489,  8.2288904,  8.2419720,  8.2550964,  8.2682619,  8.2814703,  8.2947206,  8.3080139,  8.3213501,  8.3347273,  8.3481483,  8.3616133,  8.3751221,  8.3886738,  8.4022703,  8.4159107,  8.4295940,  8.4433231,  8.4570971,  8.4709158,  8.4847803,  8.4986897,  8.5126448,  8.5266457,  8.5406923,  8.5547867,  8.5689268,  8.5831137,  8.5973482,  8.6116295,  8.6259575,  8.6403341,  8.6547585,  8.6692324,  8.6837530,  8.6983232,  8.7129421,  8.7276096,  8.7423277,  8.7570953,  8.7719135,  8.7867804,  8.8016987,  8.8166676,  8.8316870,  8.8467579,  8.8618813,  8.8770561,  8.8922825,  8.9075613,  8.9228926,  8.9382763,  8.9537134,  8.9692049,  8.9847498,  9.0003481,  9.0160007,  9.0317087,  9.0474701,  9.0632877,  9.0791597,  9.0950880,  9.1110725,  9.1271133,  9.1432114,  9.1593647,  9.1755753,  9.1918449,  9.2081718,  9.2245560,  9.2409992,  9.2575016,  9.2740612,  9.2906818,  9.3073616,  9.3241014,  9.3409014,  9.3577623,  9.3746853,  9.3916674,  9.4087124,  9.4258194,  9.4429884,  9.4602203,  9.4775152,  9.4948730,  9.5122938,  9.5297794,  9.5473309,  9.5649452,  9.5826263,  9.6003714,  9.6181831,  9.6360598,  9.6540041,  9.6720152,  9.6900940,  9.7082405,  9.7264557,  9.7447386,  9.7630892,  9.7815113,  9.8000011,  9.8185616,  9.8371925,  9.8558950,  9.8746681,  9.8935127,  9.9124298,  9.9314175,  9.9504805,  9.9696159,  9.9888258, 10.0081091, 10.0274677, 10.0469007, 10.0664082, 10.0859928, 10.1056547, 10.1253910, 10.1452065, 10.1650991, 10.1850710, 10.2051182, 10.2252474, 10.2454548, 10.2657442, 10.2861118, 10.3065615, 10.3270922, 10.3477049, 10.3684015, 10.3891792, 10.4100418, 10.4309864, 10.4520168, 10.4731321, 10.4943323, 10.5156193, 10.5369930, 10.5584545, 10.5800018, 10.6016369, 10.6233616, 10.6451750, 10.6670790, 10.6890736, 10.7111588, 10.7333345, 10.7556019, 10.7779636, 10.8004179, 10.8229656, 10.8456078, 10.8683443, 10.8911772, 10.9141064, 10.9371319, 10.9602547, 10.9834757, 11.0067949, 11.0302143, 11.0537329, 11.0773525, 11.1010714, 11.1248941, 11.1488180, 11.1728468, 11.1969786, 11.2212133, 11.2455549, 11.2700005, 11.2945538, 11.3192158, 11.3439837, 11.3688612, 11.3938465, 11.4189434, 11.4441509, 11.4694700, 11.4949017, 11.5204458, 11.5461044, 11.5718765, 11.5977631, 11.6237688, 11.6498880, 11.6761274, 11.7024851, 11.7289610, 11.7555561, 11.7822733, 11.8091135, 11.8360748, 11.8631592, 11.8903685, 11.9177027, 11.9451618, 11.9727488, 12.0004635, 12.0283079, 12.0562801, 12.0843830, 12.1126184,  
12.5, 12.7, 12.8, 13.2, 13.5, 13.9, 14.3, 14.7, 14.9, 15.4, 
15.9, 16.1, 16.7, 16.9, 17.2, 17.5, 17.9, 18.2, 18.5, 18.9, 
19.6, 20.0, 20.4, 20.8, 21.3, 22.2, 22.7, 23.3, 24.4, 25.0  ;

 bnd_PaW75 =
 25.000, 24.390, 23.256, 22.727, 22.222, 21.277, 20.833, 20.408, 20.000, 19.608, 18.868, 18.519, 18.182, 17.857, 17.544, 17.241, 16.949, 16.667, 16.129, 15.873, 15.385, 14.925, 14.706, 14.286, 13.889, 13.514, 13.158, 12.821, 12.658, 12.500, 12.195, 11.905, 11.765, 11.494, 11.442, 11.364, 11.236, 11.111, 10.989, 10.870, 10.753, 10.638, 10.526, 10.417, 10.384, 10.309, 10.204, 10.101,  9.901,  9.804,  9.709,  9.615,  9.524,  9.434,  9.346,  9.259,  9.174,  9.091,  9.009,  8.929,  8.850,  8.696,  8.621,  8.547,  8.403,  8.264,  8.130,  8.065,  8.000,  7.874,  7.752,7.634,  7.576,  7.463,  7.353,  7.299,  7.194,  7.092,  6.993,  6.897,  6.803,  6.711,  6.667,  6.623,  6.579,  6.536,  6.494,  6.410,  6.329,  6.250,  6.211,  6.173,  6.135,  6.098,  6.061,  6.024,  5.952,  5.882,  5.814,  5.747,  5.682,  5.650,  5.618,  5.556,  5.495,  5.435,  5.376,  5.319,  5.263,  5.181,  5.102,  4.950,  4.808,  4.717,  4.587,  4.464,  4.367,  4.292,  4.274,  4.219,  4.149,  4.082,  4.000,  3.953,  3.906,  3.861,  3.846,  3.817,3.759,  3.690,  3.623,  3.559,  3.472,  3.413,  3.344,  3.279,  3.175,  3.077,  3.021,  2.985,  2.941,  2.915,  2.882,  2.841,  2.833,  2.770,  2.762,  2.725,  2.688,  2.632,  2.564,  2.500,  2.439,  2.381,  2.326,  2.273,  2.222,  2.174,  2.128,  
2.083,  2.041,  2.000,  1.961,  1.923,  1.887,  1.852,  1.818,  
1.786,  1.754,  1.724,  1.695,  1.667,  1.639,  1.613,  1.587,  1.562,  1.538,  
1.515,  1.493,  1.471,  1.449,  1.429,  1.408,  1.389,  1.370,  1.351,  1.333,  
1.316,  1.299,  1.282,  1.266,  1.250,  1.220,  1.190,  1.163,  1.136,  1.111,  
1.087,  1.064,  1.042,  1.020,  1.000,   .980,   .962,   .943,   .926,   .909,   
 .893,   .877,   .862,   .847,   .833,   .820,   .806,   .794,   .781,   .769,   
 .758,   .746,   .735,   .725,   .714,   .702,   .556,   .449,   .445,   .360  ;
 
 bnd_HSL88 =
 0.200, 0.250, 0.300, 0.337, 0.400, 0.488, 0.515, 0.550, 0.633, 0.694, 0.860, 1.060, 
 1.300, 1.536, 1.800, 2.000, 2.250, 2.500, 2.700, 3.000, 3.200, 3.392, 3.500, 3.750, 
 4.000, 4.500, 5.000, 5.500, 6.000, 6.200, 6.500, 7.200, 7.900, 8.200, 8.500, 8.700, 
 9.000, 9.200, 9.500, 9.800,10.000,10.591,11.000,11.500,12.500,13.000,14.000,14.800,
15.000,16.400,17.200,18.000,18.500,20.000,21.300,22.500,25.000  ;

 idx_rfr_H2SO4_210K_61_NNM98_img = 
1.07e-8, 1.07e-8, 1.07e-8, 1.07e-8,
0.00E+00,  0.00E+00,  0.00E+00,  0.00E+00,  2.07E-08,  2.79E-08,  3.58E-08,  4.80E-08,  6.83E-08,  7.84E-08,  
8.20E-08,  8.39E-08,  8.46E-08,  8.79E-08,  9.98E-08,  1.24E-07,  1.58E-07,  1.83E-07,  2.02E-07,  2.33E-07,  
2.84E-07,  3.62E-07,  6.05E-07,  1.03E-06,  1.41E-06,  1.53E-06,  1.52E-06,  1.48E-06,  1.50E-06,  1.60E-06,  
1.84E-06,  2.46E-06,  4.05E-06,  4.95E-06,  5.63E-06,  6.94E-06,  7.75E-06,  8.93E-06,  1.05E-05,  1.27E-05,  
1.59E-05,  1.98E-05,  2.59E-05,  3.89E-05,  6.16E-05,  8.78E-05,  1.02E-04,  1.10E-04,  1.17E-04,  1.25E-04,  
1.38E-04,  1.55E-04,  1.76E-04,  2.02E-04,  2.34E-04,  2.72E-04,  3.14E-04,  3.61E-04,  4.24E-04,  4.86E-04,  
5.37E-04,  5.95E-04,  7.96E-04,  1.11E-03,  1.24E-03,  1.26E-03,  1.30E-03,  1.35E-03,
 0.00194,  0.00190,  0.00164,  0.00141,  0.00187,  0.00205,  0.00153,  0.00128,  0.00130,  0.00117,  0.00133,  0.00181,  0.00183,  0.00183,  0.00203,  0.00175,  0.00162,  0.00182,  0.00167,  0.00171,  0.00196,  0.00155,  0.00113,  0.00161,  0.00274,  0.00298,  0.00214,  0.00159,  0.00188,  0.00183,  0.00128,  0.00059,  0.00038,  0.00119,  0.00220,  0.00256,  0.00240,  0.00201,  0.00180,  0.00200,  0.00205,  0.00175,  0.00151,  0.00153,  0.00190,  0.00242,  0.00282,  0.00287,  0.00300,  0.00265,  0.00212,  0.00203,  0.00201,  0.00187,  0.00196,  0.00243,  0.00252,  0.00238,  0.00245,  0.00238,  0.00233,  0.00218,  0.00184,  0.00145,  0.00097,  0.00057,  0.00024,  0.00039,  0.00163,  0.00229,  0.00186,  0.00115,  0.00093,  0.00144,  0.00167,  0.00141,  0.00106,  0.00085,  0.00119,  0.00168,  0.00158,  0.00132,  0.00137,  0.00182,  0.00218,  0.00198,  0.00155,  0.00124,  0.00080,  0.00057,  0.00068,  0.00054,  0.00060,  0.00113,  0.00143,  0.00144,  0.00170,  0.00198,  0.00192,  0.00160,  0.00146,  0.00174,  0.00177,  0.00184,  0.00202,  0.00155,  0.00144,  0.00225,  0.00254,  0.00228,  0.00236,  0.00252,  0.00191,  0.00138,  0.00183,  0.00255,  0.00269,  0.00214,  0.00118,  0.00053,  0.00076,  0.00155,  0.00207,  0.00238,  0.00262,  0.00233,  0.00197,  0.00216,  0.00219,  0.00163,  0.00100,  0.00128,  0.00167,  0.00132,  0.00052,  0.00006,  0.00017,  0.00035,  0.00008,  0.00026,  0.00133,  0.00150,  0.00139,  0.00163,  0.00142,  0.00107,  0.00115,  0.00145,  0.00186,  0.00208,  0.00182,  0.00156,  0.00132,  0.00112,  0.00148,  0.00220,  0.00238,  0.00185,  0.00090,  0.00052,  0.00179,  0.00293,  0.00256,  0.00175,  0.00180,  0.00251,  0.00299,  0.00300,  0.00302,  0.00320,  0.00296,  0.00241,  0.00230,  0.00219,  0.00188,  0.00172,  0.00221,  0.00239,  0.00167,  0.00177,  0.00271,  0.00279,  0.00235,  0.00221,  0.00229,  0.00205,  0.00181,  0.00176,  0.00196,  0.00233,  0.00230,  0.00200,  0.00130,  0.00029,  0.00062,  0.00219,  0.00260,  0.00208,  0.00207,  0.00250,  0.00246,  0.00216,  0.00182,  0.00144,  0.00127,  0.00104,  0.00058,  0.00036,  0.00058,  0.00094,  0.00155,  0.00234,  0.00250,  0.00220,  0.00177,  0.00122,  0.00099,  0.00129,  0.00145,  0.00103,  0.00083,  0.00144,  0.00211,  0.00208,  0.00161,  0.00115,  0.00105,  0.00114,  0.00082,  0.00065,  0.00117,  0.00200,  0.00249,  0.00230,  0.00203,  0.00200,  0.00181,  0.00172,  0.00196,  0.00215,  0.00209,  0.00255,  0.00336,  0.00334,  0.00310,  0.00293,  0.00279,  0.00256,  0.00226,  0.00184,  0.00143,  0.00098,  0.00038,  0.00004,  0.00045,  0.00140,  0.00219,  0.00223,  0.00173,  0.00139,  0.00132,  0.00121,  0.00104,  0.00092,  0.00110,  0.00171,  0.00216,  0.00232,  0.00225,  0.00188,  0.00160,  0.00156,  0.00118,  0.00083,  0.00102,  0.00132,  0.00196,  0.00271,  0.00255,  0.00200,  0.00183,  0.00181,  0.00181,  0.00233,  0.00315,  0.00320,  0.00278,  0.00213,  0.00148,  0.00145,  0.00165,  0.00165,  0.00199,  0.00256,  0.00252,  0.00185,  0.00154,  0.00172,  0.00195,  0.00214,  0.00214,  0.00136,  0.00024,  0.00072,  0.00197,  0.00212,  0.00189,  0.00182,  0.00201,  0.00224,  0.00228,  0.00243,  0.00271,  0.00266,  0.00262,  0.00287,  0.00344,  0.00418,  0.00405,  0.00343,  0.00301,  0.00298,  0.00316,  0.00309,  0.00288,  0.00275,  0.00275,  0.00293,  0.00342,  0.00384,  0.00393,  0.00390,  0.00375,  0.00364,  0.00348,  0.00300,  0.00248,  0.00253,  0.00290,  0.00272,  0.00261,  0.00318,  0.00326,  0.00283,  0.00295,  0.00319,  0.00307,  0.00354,  0.00420,  0.00384,  0.00329,  0.00295,  0.00268,  0.00226,  0.00217,  0.00254,  0.00280,  0.00298,  0.00305,  0.00294,  0.00275,  0.00268,  0.00272,  0.00264,  0.00259,  0.00302,  0.00376,  0.00389,  0.00333,  0.00297,  0.00314,  0.00351,  0.00356,  0.00314,  0.00274,  0.00300,  0.00341,  0.00361,  0.00359,  0.00321,  0.00340,  0.00414,  0.00446,  0.00415,  0.00399,  0.00402,  0.00400,  0.00386,  0.00343,  0.00312,  0.00320,  0.00365,  0.00377,  0.00350,  0.00366,  0.00395,  0.00399,  0.00374,  0.00348,  0.00351,  0.00387,  0.00428,  0.00446,  0.00441,  0.00411,  0.00384,  0.00374,  0.00379,  0.00401,  0.00417,  0.00429,  0.00435,  0.00430,  0.00414,  0.00394,  0.00405,  0.00410,  0.00394,  0.00399,  0.00378,  0.00321,  0.00298,  0.00317,  0.00321,  0.00314,  0.00327,  0.00347,  0.00355,  0.00321,  0.00278,  0.00296,  0.00337,  0.00364,  0.00390,  0.00411,  0.00419,  0.00401,  0.00395,  0.00436,  0.00478,  0.00463,  0.00426,  0.00416,  0.00395,  0.00386,  0.00416,  0.00434,  0.00441,  0.00444,  0.00415,  0.00404,  0.00417,  0.00414,  0.00419,  0.00429,  0.00448,  0.00474,  0.00479,  0.00489,  0.00479,  0.00455,  0.00446,  0.00434,  0.00427,  0.00427,  0.00442,  0.00454,  0.00447,  0.00434,  0.00408,  0.00411,  0.00417,  0.00406,  0.00401,  0.00413,  0.00405,  0.00395,  0.00406,  0.00420,  0.00426,  0.00430,  0.00447,  0.00471,  0.00493,  0.00519,  0.00497,  0.00458,  0.00483,  0.00492,  0.00455,  0.00449,  0.00457,  0.00467,  0.00475,  0.00444,  0.00439,  0.00457,  0.00455,  0.00438,  0.00397,  0.00384,  0.00407,  0.00433,  0.00427,  0.00418,  0.00437,  0.00449,  0.00437,  0.00442,  0.00466,  0.00485,  0.00483,  0.00503,  0.00503,  0.00466,  0.00463,  0.00470,  0.00472,  0.00479,  0.00471,  0.00450,  0.00460,  0.00489,  0.00485,  0.00480,  0.00487,  0.00497,  0.00501,  0.00505,  0.00519,  0.00540,  0.00578,  0.00594,  0.00607,  0.00627,  0.00627,  0.00629,  0.00632,  0.00666,  0.00708,  0.00756,  0.00793,  0.00796,  0.00817,  0.00872,  0.00914,  0.00960,  0.01040,  0.01082,  0.01146,  0.01225,  0.01277,  0.01371,  0.01471,  0.01554,  0.01670,  0.01772,  0.01860,  0.01963,  0.02103,  0.02265,  0.02372,  0.02454,  0.02526,  0.02626,  0.02748,  0.02879,  0.03008,  0.03121,  0.03245,  0.03333,  0.03470,  0.03646,  0.03775,  0.03877,  0.03992,  0.04150,  0.04303,  0.04421,  0.04522,  0.04662,  0.04803,  0.04951,  0.05110,  0.05238,  0.05404,  0.05558,  0.05673,  0.05807,  0.05947,  0.06070,  0.06189,  0.06341,  0.06532,  0.06689,  0.06834,  0.06973,  0.07070,  0.07207,  0.07370,  0.07526,  0.07679,  0.07817,  0.07912,  0.08041,  0.08237,  0.08388,  0.08554,  0.08718,  0.08843,  0.08980,  0.09137,  0.09288,  0.09373,  0.09504,  0.09710,  0.09886,  0.10031,  0.10185,  0.10332,  0.10485,  0.10649,  0.10760,  0.10849,  0.11021,  0.11176,  0.11296,  0.11437,  0.11588,  0.11748,  0.11857,  0.12033,  0.12187,  0.12317,  0.12501,  0.12604,  0.12737,  0.12932,  0.13111,  0.13261,  0.13327,  0.13401,  0.13562,  0.13728,  0.13886,  0.14012,  0.14104,  0.14240,  0.14408,  0.14580,  0.14666,  0.14765,  0.14922,  0.15036,  0.15196,  0.15288,  0.15326,  0.15482,  0.15685,  0.15836,  0.15942,  0.16042,  0.16149,  0.16235,  0.16339,  0.16462,  0.16546,  0.16635,  0.16727,  0.16858,  0.16963,  0.17040,  0.17148,  0.17268,  0.17423,  0.17477,  0.17512,  0.17632,  0.17689,  0.17723,  0.17861,  0.17932,  0.18006,  0.18081,  0.18150,  0.18219,  0.18281,  0.18342,  0.18398,  0.18455,  0.18511,  0.18567,  0.18621,  0.18673,  0.18720,  0.18764,  0.18808,  0.18848,  0.18884,  0.18918,  0.18952,  0.18985,  0.19014,  0.19043,  0.19071,  0.19101,  0.19128,  0.19152,  0.19175,  0.19198,  0.19219,  0.19241,  0.19260,  0.19277,  0.19290,  0.19305,  0.19319,  0.19336,  0.19355,  0.19373,  0.19388,  0.19402,  0.19415,  0.19427,  0.19438,  0.19450,  0.19461,  0.19472,  0.19484,  0.19495,  0.19505,  0.19517,  0.19527,  0.19536,  0.19545,  0.19556,  0.19567,  0.19581,  0.19593,  0.19601,  0.19609,  0.19617,  0.19624,  0.19630,  0.19637,  0.19643,  0.19647,  0.19652,  0.19655,  0.19658,  0.19660,  0.19660,  0.19657,  0.19651,  0.19644,  0.19638,  0.19632,  0.19628,  0.19625,  0.19623,  0.19620,  0.19615,  0.19611,  0.19606,  0.19601,  0.19595,  0.19588,  0.19582,  0.19574,  0.19564,  0.19554,  0.19545,  0.19533,  0.19523,  0.19514,  0.19503,  0.19494,  0.19484,  0.19469,  0.19453,  0.19438,  0.19425,  0.19412,  0.19399,  0.19386,  0.19375,  0.19361,  0.19348,  0.19335,  0.19322,  0.19311,  0.19300,  0.19287,  0.19275,  0.19264,  0.19252,  0.19240,  0.19228,  0.19213,  0.19201,  0.19192,  0.19180,  0.19167,  0.19154,  0.19140,  0.19126,  0.19112,  0.19097,  0.19081,  0.19066,  0.19053,  0.19041,  0.19028,  0.19017,  0.19006,  0.18997,  0.18990,  0.18983,  0.18975,  0.18966,  0.18956,  0.18949,  0.18942,  0.18933,  0.18926,  0.18920,  0.18914,  0.18908,  0.18902,  0.18896,  0.18891,  0.18888,  0.18883,  0.18880,  0.18878,  0.18875,  0.18873,  0.18871,  0.18869,  0.18868,  0.18866,  0.18867,  0.18867,  0.18867,  0.18870,  0.18873,  0.18875,  0.18877,  0.18878,  0.18879,  0.18880,  0.18881,  0.18883,  0.18886,  0.18886,  0.18886,  0.18885,  0.18882,  0.18879,  0.18877,  0.18875,  0.18873,  0.18870,  0.18868,  0.18865,  0.18861,  0.18855,  0.18847,  0.18837,  0.18826,  0.18815,  0.18801,  0.18784,  0.18767,  0.18750,  0.18732,  0.18712,  0.18692,  0.18670,  0.18652,  0.18638,  0.18626,  0.18613,  0.18600,  0.18592,  0.18585,  0.18579,  0.18571,  0.18561,  0.18553,  0.18548,  0.18546,  0.18543,  0.18540,  0.18541,  0.18545,  0.18551,  0.18561,  0.18576,  0.18591,  0.18613,  0.18638,  0.18667,  0.18700,  0.18733,  0.18767,  0.18802,  0.18840,  0.18881,  0.18923,  0.18966,  0.19008,  0.19051,  0.19093,  0.19136,  0.19179,  0.19221,  0.19262,  0.19302,  0.19341,  0.19379,  0.19417,  0.19455,  0.19490,  0.19521,  0.19549,  0.19576,  0.19600,  0.19622,  0.19644,  0.19665,  0.19683,  0.19701,  0.19720,  0.19739,  0.19757,  0.19776,  0.19798,  0.19820,  0.19842,  0.19864,  0.19883,  0.19899,  0.19915,  0.19928,  0.19940,  0.19948,  0.19955,  0.19962,  0.19971,  0.19980,  0.19989,  0.19999,  0.20010,  0.20023,  0.20034,  0.20043,  0.20053,  0.20063,  0.20072,  0.20084,  0.20094,  0.20104,  0.20111,  0.20116,  0.20122,  0.20124,  0.20122,  0.20120,  0.20118,  0.20114,  0.20107,  0.20099,  0.20088,  0.20075,  0.20057,  0.20036,  0.20014,  0.19994,  0.19974,  0.19954,  0.19934,  0.19912,  0.19885,  0.19859,  0.19833,  0.19806,  0.19779,  0.19752,  0.19725,  0.19698,  0.19671,  0.19644,  0.19615,  0.19586,  0.19555,  0.19526,  0.19495,  0.19462,  0.19430,  0.19396,  0.19364,  0.19331,  0.19298,  0.19263,  0.19228,  0.19192,  0.19157,  0.19121,  0.19083,  0.19047,  0.19012,  0.18976,  0.18939,  0.18900,  0.18863,  0.18828,  0.18794,  0.18761,  0.18729,  0.18697,  0.18663,  0.18629,  0.18595,  0.18561,  0.18527,  0.18494,  0.18463,  0.18432,  0.18400,  0.18367,  0.18333,  0.18300,  0.18267,  0.18235,  0.18207,  0.18179,  0.18150,  0.18123,  0.18094,  0.18067,  0.18040,  0.18011,  0.17983,  0.17957,  0.17932,  0.17905,  0.17880,  0.17855,  0.17831,  0.17807,  0.17784,  0.17761,  0.17739,  0.17717,  0.17696,  0.17676,  0.17656,  0.17637,  0.17619,  0.17601,  0.17585,  0.17567,  0.17549,  0.17531,  0.17512,  0.17496,  0.17479,  0.17462,  0.17446,  0.17432,  0.17419,  0.17407,  0.17395,  0.17381,  0.17369,  0.17357,  0.17343,  0.17329,  0.17315,  0.17299,  0.17285,  0.17272,  0.17258,  0.17243,  0.17230,  0.17216,  0.17202,  0.17184,  0.17167,  0.17151,  0.17136,  0.17121,  0.17105,  0.17088,  0.17072,  0.17055,  0.17038,  0.17022,  0.17005,  0.16990,  0.16974,  0.16957,  0.16940,  0.16924,  0.16908,  0.16893,  0.16878,  0.16861,  0.16843,  0.16828,  0.16790,  0.16764,  0.16758,  0.16763,  0.16741,  0.16707,  0.16702,  0.16714,  0.16717,  0.16679,  0.16669,  0.16676,  0.16654,  0.16659,  0.16649,  0.16608,  0.16566,  0.16557,  0.16571,  0.16541,  0.16506,  0.16509,  0.16506,  0.16480,  0.16442,  0.16396,  0.16398,  0.16438,  0.16439,  0.16441,  0.16461,  0.16431,  0.16397,  0.16392,  0.16389,  0.16396,  0.16413,  0.16393,  0.16367,  0.16344,  0.16336,  0.16361,  0.16318,  0.16256,  0.16245,  0.16220,  0.16210,  0.16220,  0.16188,  0.16154,  0.16140,  0.16133,  0.16119,  0.16104,  0.16104,  0.16100,  0.16082,  0.16083,  0.16073,  0.16037,  0.16033,  0.16017,  0.15995,  0.15974,  0.15942,  0.15928,  0.15922,  0.15894,  0.15872,  0.15881,  0.15885,  0.15875,  0.15867,  0.15857,  0.15836,  0.15806,  0.15806,  0.15835,  0.15830,  0.15843,  0.15892,  0.15880,  0.15854,  0.15864,  0.15836,  0.15808,  0.15804,  0.15796,  0.15807,  0.15819,  0.15828,  0.15829,  0.15862,  0.15887,  0.15869,  0.15863,  0.15849,  0.15847,  0.15875,  0.15895,  0.15914,  0.15953,  0.15972,  0.15974,  0.15960,  0.15939,  0.15952,  0.15980,  0.16011,  0.16040,  0.16078,  0.16092,  0.16108,  0.16156,  0.16156,  0.16103,  0.16084,  0.16101,  0.16126,  0.16169,  0.16201,  0.16221,  0.16232,  0.16255,  0.16259,  0.16231,  0.16268,  0.16318,  0.16324,  0.16361,  0.16387,  0.16369,  0.16377,  0.16402,  0.16426,  0.16441,  0.16444,  0.16471,  0.16521,  0.16524,  0.16510,  0.16518,  0.16539,  0.16560,  0.16579,  0.16611,  0.16626,  0.16644,  0.16646,  0.16633,  0.16665,  0.16646,  0.16639,  0.16699,  0.16705,  0.16689,  0.16704,  0.16714,  0.16708,  0.16725,  0.16741,  0.16730,  0.16739,  0.16778,  0.16785,  0.16767,  0.16725,  0.16717,  0.16784,  0.16809,  0.16799,  0.16795,  0.16789,  0.16806,  0.16819,  0.16812,  0.16795,  0.16792,  0.16797,  0.16780,  0.16785,  0.16790,  0.16781,  0.16773,  0.16776,  0.16789,  0.16783,  0.16784,  0.16765,  0.16744,  0.16715,  0.16667,  0.16693,  0.16710,  0.16667,  0.16663,  0.16644,  0.16595,  0.16584,  0.16582,  0.16575,  0.16543,  0.16492,  0.16471,  0.16453,  0.16416,  0.16415,  0.16414,  0.16398,  0.16376,  0.16340,  0.16339,  0.16329,  0.16313,  0.16281,  0.16239,  0.16226,  0.16210,  0.16211,  0.16230,  0.16216,  0.16191,  0.16163,  0.16127,  0.16118,  0.16129,  0.16131,  0.16102,  0.16096,  0.16086,  0.16071,  0.16075,  0.16061,  0.16060,  0.16047,  0.16029,  0.16012,  0.15990,  0.15983,  0.16004,  0.16016,  0.16010,  0.16020,  0.16008,  0.15987,  0.15979,  0.15970,  0.15962,  0.15953,  0.15949,  0.15939,  0.15943,  0.15973,  0.15965,  0.15944,  0.15950,  0.15960,  0.15980,  0.15990,  0.15993,  0.15988,  0.16017,  0.16060,  0.16056,  0.16052,  0.16074,  0.16111,  0.16134,  0.16149,  0.16171,  0.16179,  0.16172,  0.16185,  0.16211,  0.16243,  0.16282,  0.16300,  0.16328,  0.16373,  0.16382,  0.16399,  0.16443,  0.16458,  0.16484,  0.16538,  0.16584,  0.16616,  0.16642,  0.16676,  0.16721,  0.16783,  0.16814,  0.16836,  0.16876,  0.16922,  0.16987,  0.17036,  0.17076,  0.17141,  0.17208,  0.17249,  0.17285,  0.17334,  0.17412,  0.17496,  0.17554,  0.17609,  0.17667,  0.17716,  0.17769,  0.17849,  0.17949,  0.18021,  0.18092,  0.18182,  0.18253,  0.18325,  0.18410,  0.18497,  0.18580,  0.18673,  0.18772,  0.18863,  0.18953,  0.19052,  0.19136,  0.19242,  0.19360,  0.19457,  0.19575,  0.19700,  0.19818,  0.19922,  0.20018,  0.20134,  0.20286,  0.20429,  0.20539,  0.20646,  0.20797,  0.20986,  0.21098,  0.21174,  0.21328,  0.21469,  0.21598,  0.21773,  0.21908,  0.22041,  0.22210,  0.22366,  0.22516,  0.22677,  0.22835,  0.22987,  0.23157,  0.23295,  0.23435,  0.23608,  0.23794,  0.23982,  0.24140,  0.24315,  0.24489,  0.24616,  0.24784,  0.25000,  0.25200,  0.25379,  0.25567,  0.25751,  0.25902,  0.26074,  0.26257,  0.26434,  0.26621,  0.26813,  0.27005,  0.27201,  0.27384,  0.27559,  0.27751,  0.27920,  0.28099,  0.28273,  0.28429,  0.28614,  0.28836,  0.29041,  0.29211,  0.29393,  0.29613,  0.29813,  0.29959,  0.30172,  0.30394,  0.30550,  0.30718,  0.30914,  0.31107,  0.31305,  0.31509,  0.31703,  0.31879,  0.32042,  0.32188,  0.32329,  0.32508,  0.32685,  0.32847,  0.33005,  0.33183,  0.33365,  0.33533,  0.33693,  0.33832,  0.33922,  0.33975,  0.34097,  0.34246,  0.34360,  0.34476,  0.34560,  0.34653,  0.34764,  0.34784,  0.34834,  0.34973,  0.35052,  0.35108,  0.35182,  0.35200,  0.35192,  0.35227,  0.35274,  0.35299,  0.35250,  0.35146,  0.35106,  0.35065,  0.34957,  0.34858,  0.34779,  0.34688,  0.34581,  0.34431,  0.34267,  0.34099,  0.33894,  0.33670,  0.33448,  0.33235,  0.33074,  0.32864,  0.32577,  0.32347,  0.32079,  0.31808,  0.31544,  0.31249,  0.30995,  0.30734,  0.30438,  0.30133,  0.29833,  0.29511,  0.29211,  0.28937,  0.28688,  0.28445,  0.28108,  0.27712,  0.27425,  0.27160,  0.26843,  0.26542,  0.26229,  0.25947,  0.25650,  0.25324,  0.25052,  0.24780,  0.24452,  0.24165,  0.23899,  0.23577,  0.23268,  0.23015,  0.22761,  0.22434,  0.22154,  0.21871,  0.21566,  0.21345,  0.21137,  0.20946,  0.20739,  0.20493,  0.20280,  0.20090,  0.19910,  0.19737,  0.19565,  0.19408,  0.19265,  0.19150,  0.19045,  0.18935,  0.18852,  0.18798,  0.18714,  0.18630,  0.18599,  0.18525,  0.18433,  0.18319,  0.18267,  0.18339,  0.18288,  0.18198,  0.18208,  0.18165,  0.18121,  0.18143,  0.18158,  0.18163,  0.18158,  0.18186,  0.18204,  0.18132,  0.18098,  0.18124,  0.18142,  0.18186,  0.18220,  0.18240,  0.18315,  0.18398,  0.18416,  0.18444,  0.18513,  0.18549,  0.18590,  0.18666,  0.18741,  0.18814,  0.18861,  0.18898,  0.18962,  0.19032,  0.19093,  0.19148,  0.19228,  0.19302,  0.19347,  0.19406,  0.19464,  0.19527,  0.19589,  0.19622,  0.19678,  0.19757,  0.19847,  0.19925,  0.19990,  0.20064,  0.20156,  0.20240,  0.20287,  0.20346,  0.20432,  0.20493,  0.20522,  0.20592,  0.20688,  0.20794,  0.20885,  0.20951,  0.21023,  0.21097,  0.21181,  0.21309,  0.21452,  0.21525,  0.21536,  0.21529,  0.21599,  0.21750,  0.21855,  0.21966,  0.22110,  0.22184,  0.22199,  0.22285,  0.22437,  0.22532,  0.22638,  0.22772,  0.22876,  0.23012,  0.23225,  0.23459,  0.23651,  0.23826,  0.24017,  0.24162,  0.24309,  0.24475,  0.24631,  0.24832,  0.25033,  0.25251,  0.25488,  0.25683,  0.25815,  0.25950,  0.26045,  0.26207,  0.26547,  0.26871,  0.27194,  0.27506,  0.27672,  0.27743,  0.27807,  0.27889,  0.28007,  0.28130,  0.28280,  0.28486,  0.28721,  0.29045,  0.29354,  0.29575,  0.29831,  0.30099,  0.30363,  0.30643,  0.30891,  0.31112,  0.31367,  0.31570,  0.31749,  0.31983,  0.32183,  0.32321,  0.32431,  0.32548,  0.32698,  0.32855,  0.32959,  0.33057,  0.33165,  0.33282,  0.33395,  0.33469,  0.33571,  0.33759,  0.33908,  0.33990,  0.34143,  0.34310,  0.34469,  0.34695,  0.34939,  0.35210,  0.35542,  0.35916,  0.36352,  0.36854,  0.37439,  0.37972,  0.38600,  0.39376,  0.40047,  0.40731,  0.41425,  0.42247,  0.43220,  0.44128,  0.45128,  0.46228,  0.47310,  0.48360,  0.49441,  0.50536,  0.51665,  0.52818,  0.53957,  0.55079,  0.56184,  0.57265,  0.58325,  0.59359,  0.60376,  0.61364,  0.62302,  0.63210,  0.64112,  0.65020,  0.65942,  0.66860,  0.67720,  0.68509,  0.69271,  0.70064,  0.70931,  0.71834,  0.72751,  0.73662,  0.74512,  0.75392,  0.76325,  0.77303,  0.78356,  0.79398,  0.80426,  0.81380,  0.82208,  0.82938,  0.83596,  0.84309,  0.85046,  0.85750,  0.86357,  0.86730,  0.86919,  0.86995,  0.86973,  0.86867,  0.86799,  0.86792,  0.86743,  0.86684,  0.86521,  0.86184,  0.85761,  0.85460,  0.85360,  0.85220,  0.85029,  0.84873,  0.84547,  0.84331,  0.84540,  0.84866,  0.85023,  0.85062,  0.85244,  0.85402,  0.85500,  0.85912,  0.86260,  0.86307,  0.86378,  0.86723,  0.87236,  0.87508,  0.87609,  0.87403,  0.86808,  0.86358,  0.86344,  0.86603,  0.86747,  0.86908,  0.87252,  0.87590,  0.88173,  0.89071,  0.90053,  0.91269,  0.92782,  0.94180,  0.95291,  0.96394,  0.97603,  0.98815,  0.99995,  1.01088,  1.01929,  1.02575,  1.03139,  1.03465,  1.03548,  1.03507,  1.03372,  1.03200,  1.02863,  1.02186,  1.01251,  1.00196,  0.98831,  0.97066,  0.95088,  0.93035,  0.90983,  0.89007,  0.87089,  0.85056,  0.82838,  0.80590,  0.78323,  0.75979,  0.73627,  0.71347,  0.69127,  0.66919,  0.64842,  0.63041,  0.61523,  0.60170,  0.58898,  0.57940,  0.57469,  0.57369,  0.57349,  0.57084,  0.56352,  0.54981,  0.53902,  0.52653,  0.51352,  0.50404,  0.49621,  0.48660,  0.47801,  0.46829,  0.45934,  0.45200,  0.44355,  0.43402,  0.42654,  0.42485,  0.42105,  0.41596,  0.41362,  0.41013,  0.40720,  0.40743,  0.40795,  0.40863,  0.40992,  0.41161,  0.41592,  0.42136,  0.42561,  0.43022,  0.43766,  0.44588,  0.45475,  0.46344,  0.47216,  0.48120,  0.48899,  0.49496,  0.50046,  0.50791,  0.51218,  0.51269,  0.51117,  0.50756,  0.50300,  0.49833,  0.49240,  0.48244,  0.47116,  0.46015,  0.44790,  0.43656,  0.42467,  0.40952,  0.39504,  0.38243,  0.37376,  0.36840,  0.36320,  0.35644,  0.34848,  0.33970,  0.33049,  0.32121,  0.31224,  0.30396,  0.29674,  0.29096,  0.28628,  0.28285,  0.28052,  0.27875,  0.27705,  0.27606,  0.27569,  0.27477,  0.27342,  0.27173,  0.26984,  0.26785,  0.26589,  
0.158,    0.157,    0.157,    0.16,     0.165,    0.171,    0.173,    0.183,    0.191,    0.221,    
0.299,    0.352,    0.479,    0.564,    0.594,    0.554,    0.457,    0.362,    0.299,    0.261,    
0.238,    0.235,    0.24,     0.257,    0.29,     0.329,    0.32,     0.3,      0.226,    0.2  ;
 
 idx_rfr_H2SO4_210K_61_NNM98_rl = 
1.526, 1.512, 1.496, 1.484,
1.452,  1.438,  1.432,  1.431,  1.428,  1.427,  1.427,  1.427,  1.427,  1.427,  
1.427,  1.427,  1.427,  1.427,  1.427,  1.426,  1.426,  1.425,  1.425,  1.425,  
1.424,  1.424,  1.423,  1.423,  1.422,  1.422,  1.421,  1.421,  1.420,  1.419,  
1.418,  1.417,  1.416,  1.416,  1.415,  1.413,  1.413,  1.412,  1.411,  1.411,  
1.410,  1.410,  1.409,  1.408,  1.407,  1.406,  1.406,  1.405,  1.404,  1.403,  
1.403,  1.402,  1.400,  1.399,  1.398,  1.398,  1.397,  1.396,  1.394,  1.393,  
1.392,  1.391,  1.389,  1.388,  1.386,  1.384,  1.382,  1.380, 
 1.38800,  1.38781,  1.38759,  1.38716,  1.38688,  1.38713,  1.38720,  1.38688,  1.38656,  1.38623,  1.38581,  1.38571,  1.38578,  1.38576,  1.38582,  1.38586,  1.38563,  1.38552,  1.38543,  1.38526,  1.38533,  1.38539,  1.38482,  1.38408,  1.38421,  1.38511,  1.38556,  1.38519,  1.38493,  1.38514,  1.38523,  1.38473,  1.38370,  1.38288,  1.38290,  1.38345,  1.38390,  1.38396,  1.38370,  1.38353,  1.38362,  1.38362,  1.38330,  1.38282,  1.38242,  1.38235,  1.38257,  1.38286,  1.38322,  1.38353,  1.38346,  1.38317,  1.38301,  1.38278,  1.38244,  1.38239,  1.38260,  1.38270,  1.38272,  1.38281,  1.38293,  1.38309,  1.38320,  1.38318,  1.38297,  1.38257,  1.38184,  1.38086,  1.38051,  1.38114,  1.38181,  1.38169,  1.38109,  1.38076,  1.38095,  1.38113,  1.38096,  1.38046,  1.38003,  1.38007,  1.38028,  1.38014,  1.37977,  1.37963,  1.37993,  1.38034,  1.38046,  1.38039,  1.38013,  1.37968,  1.37931,  1.37896,  1.37844,  1.37813,  1.37814,  1.37809,  1.37799,  1.37812,  1.37836,  1.37833,  1.37802,  1.37782,  1.37776,  1.37771,  1.37783,  1.37774,  1.37716,  1.37692,  1.37727,  1.37745,  1.37742,  1.37771,  1.37787,  1.37733,  1.37671,  1.37681,  1.37746,  1.37799,  1.37789,  1.37705,  1.37606,  1.37561,  1.37566,  1.37588,  1.37626,  1.37657,  1.37648,  1.37639,  1.37669,  1.37687,  1.37642,  1.37592,  1.37606,  1.37646,  1.37633,  1.37567,  1.37503,  1.37475,  1.37429,  1.37352,  1.37331,  1.37362,  1.37369,  1.37373,  1.37384,  1.37360,  1.37314,  1.37283,  1.37283,  1.37310,  1.37330,  1.37325,  1.37301,  1.37252,  1.37199,  1.37202,  1.37256,  1.37300,  1.37262,  1.37139,  1.37056,  1.37109,  1.37188,  1.37171,  1.37097,  1.37064,  1.37089,  1.37117,  1.37127,  1.37153,  1.37187,  1.37186,  1.37164,  1.37155,  1.37135,  1.37085,  1.37062,  1.37088,  1.37072,  1.37001,  1.36991,  1.37041,  1.37059,  1.37040,  1.37036,  1.37035,  1.37015,  1.36979,  1.36951,  1.36956,  1.36986,  1.37016,  1.37018,  1.36928,  1.36790,  1.36759,  1.36830,  1.36856,  1.36828,  1.36830,  1.36864,  1.36884,  1.36885,  1.36868,  1.36845,  1.36830,  1.36793,  1.36725,  1.36657,  1.36603,  1.36571,  1.36591,  1.36648,  1.36690,  1.36701,  1.36676,  1.36620,  1.36583,  1.36587,  1.36574,  1.36509,  1.36457,  1.36474,  1.36523,  1.36541,  1.36513,  1.36470,  1.36448,  1.36420,  1.36350,  1.36278,  1.36264,  1.36304,  1.36339,  1.36337,  1.36325,  1.36307,  1.36272,  1.36241,  1.36230,  1.36200,  1.36167,  1.36189,  1.36245,  1.36273,  1.36281,  1.36291,  1.36302,  1.36308,  1.36304,  1.36289,  1.36265,  1.36213,  1.36115,  1.36012,  1.35965,  1.35996,  1.36053,  1.36072,  1.36048,  1.36018,  1.35995,  1.35965,  1.35915,  1.35855,  1.35823,  1.35832,  1.35859,  1.35884,  1.35889,  1.35869,  1.35852,  1.35831,  1.35774,  1.35706,  1.35649,  1.35619,  1.35648,  1.35700,  1.35701,  1.35665,  1.35628,  1.35578,  1.35536,  1.35555,  1.35618,  1.35663,  1.35665,  1.35616,  1.35551,  1.35509,  1.35472,  1.35436,  1.35445,  1.35488,  1.35490,  1.35438,  1.35389,  1.35368,  1.35370,  1.35402,  1.35413,  1.35316,  1.35180,  1.35147,  1.35181,  1.35180,  1.35143,  1.35108,  1.35089,  1.35071,  1.35047,  1.35038,  1.35029,  1.34998,  1.34953,  1.34931,  1.34967,  1.35032,  1.35052,  1.35018,  1.34977,  1.34958,  1.34954,  1.34936,  1.34901,  1.34857,  1.34810,  1.34784,  1.34793,  1.34814,  1.34828,  1.34833,  1.34834,  1.34841,  1.34834,  1.34784,  1.34719,  1.34694,  1.34678,  1.34629,  1.34603,  1.34617,  1.34599,  1.34555,  1.34534,  1.34503,  1.34471,  1.34502,  1.34553,  1.34556,  1.34530,  1.34503,  1.34455,  1.34385,  1.34331,  1.34308,  1.34298,  1.34293,  1.34285,  1.34261,  1.34226,  1.34195,  1.34162,  1.34106,  1.34051,  1.34051,  1.34095,  1.34105,  1.34058,  1.34003,  1.33987,  1.34000,  1.33994,  1.33937,  1.33872,  1.33841,  1.33839,  1.33839,  1.33802,  1.33735,  1.33712,  1.33742,  1.33758,  1.33739,  1.33719,  1.33712,  1.33711,  1.33690,  1.33634,  1.33568,  1.33536,  1.33532,  1.33508,  1.33465,  1.33446,  1.33449,  1.33437,  1.33396,  1.33337,  1.33292,  1.33278,  1.33287,  1.33297,  1.33290,  1.33258,  1.33213,  1.33167,  1.33133,  1.33113,  1.33099,  1.33091,  1.33084,  1.33069,  1.33036,  1.33004,  1.32989,  1.32971,  1.32956,  1.32952,  1.32918,  1.32850,  1.32794,  1.32759,  1.32717,  1.32671,  1.32642,  1.32634,  1.32615,  1.32550,  1.32468,  1.32415,  1.32383,  1.32357,  1.32341,  1.32332,  1.32308,  1.32255,  1.32211,  1.32213,  1.32226,  1.32207,  1.32171,  1.32128,  1.32069,  1.32020,  1.31993,  1.31975,  1.31961,  1.31933,  1.31882,  1.31837,  1.31799,  1.31755,  1.31709,  1.31670,  1.31645,  1.31626,  1.31612,  1.31598,  1.31570,  1.31530,  1.31490,  1.31443,  1.31393,  1.31350,  1.31325,  1.31300,  1.31260,  1.31221,  1.31166,  1.31124,  1.31081,  1.31028,  1.30981,  1.30939,  1.30883,  1.30823,  1.30775,  1.30728,  1.30675,  1.30622,  1.30576,  1.30541,  1.30528,  1.30515,  1.30461,  1.30403,  1.30378,  1.30339,  1.30275,  1.30214,  1.30168,  1.30136,  1.30089,  1.30023,  1.29968,  1.29932,  1.29893,  1.29828,  1.29736,  1.29652,  1.29598,  1.29548,  1.29477,  1.29408,  1.29354,  1.29293,  1.29215,  1.29145,  1.29092,  1.29035,  1.28982,  1.28941,  1.28880,  1.28795,  1.28718,  1.28645,  1.28577,  1.28510,  1.28422,  1.28323,  1.28244,  1.28174,  1.28088,  1.27994,  1.27906,  1.27816,  1.27718,  1.27613,  1.27508,  1.27417,  1.27333,  1.27243,  1.27153,  1.27061,  1.26952,  1.26825,  1.26694,  1.26572,  1.26465,  1.26371,  1.26261,  1.26122,  1.25987,  1.25857,  1.25719,  1.25593,  1.25469,  1.25333,  1.25204,  1.25067,  1.24922,  1.24794,  1.24666,  1.24542,  1.24434,  1.24319,  1.24182,  1.24057,  1.23976,  1.23922,  1.23854,  1.23752,  1.23634,  1.23519,  1.23423,  1.23338,  1.23258,  1.23180,  1.23082,  1.22967,  1.22888,  1.22844,  1.22778,  1.22684,  1.22598,  1.22548,  1.22504,  1.22432,  1.22349,  1.22275,  1.22209,  1.22157,  1.22102,  1.22051,  1.22025,  1.21994,  1.21947,  1.21907,  1.21868,  1.21806,  1.21734,  1.21694,  1.21682,  1.21674,  1.21668,  1.21640,  1.21586,  1.21547,  1.21528,  1.21521,  1.21525,  1.21501,  1.21440,  1.21403,  1.21394,  1.21388,  1.21398,  1.21408,  1.21396,  1.21394,  1.21417,  1.21413,  1.21360,  1.21334,  1.21358,  1.21382,  1.21398,  1.21415,  1.21434,  1.21478,  1.21524,  1.21521,  1.21513,  1.21543,  1.21571,  1.21577,  1.21594,  1.21630,  1.21647,  1.21665,  1.21702,  1.21736,  1.21783,  1.21833,  1.21844,  1.21868,  1.21947,  1.22060,  1.22144,  1.22158,  1.22161,  1.22206,  1.22283,  1.22366,  1.22419,  1.22445,  1.22495,  1.22597,  1.22692,  1.22745,  1.22801,  1.22872,  1.22966,  1.23076,  1.23117,  1.23120,  1.23191,  1.23319,  1.23440,  1.23542,  1.23641,  1.23730,  1.23809,  1.23905,  1.24008,  1.24092,  1.24161,  1.24249,  1.24356,  1.24453,  1.24527,  1.24615,  1.24754,  1.24908,  1.25003,  1.25104,  1.25225,  1.25302,  1.25388,  1.25510,  1.25624,  1.25732,  1.25846,  1.25957,  1.26072,  1.26183,  1.26293,  1.26400,  1.26509,  1.26616,  1.26726,  1.26836,  1.26948,  1.27057,  1.27167,  1.27276,  1.27384,  1.27489,  1.27594,  1.27698,  1.27800,  1.27899,  1.27997,  1.28095,  1.28195,  1.28292,  1.28388,  1.28482,  1.28576,  1.28669,  1.28763,  1.28855,  1.28946,  1.29032,  1.29115,  1.29197,  1.29280,  1.29365,  1.29450,  1.29534,  1.29617,  1.29699,  1.29779,  1.29858,  1.29936,  1.30013,  1.30091,  1.30167,  1.30243,  1.30318,  1.30393,  1.30467,  1.30539,  1.30611,  1.30683,  1.30756,  1.30832,  1.30907,  1.30981,  1.31055,  1.31130,  1.31202,  1.31275,  1.31348,  1.31421,  1.31494,  1.31567,  1.31639,  1.31712,  1.31786,  1.31860,  1.31930,  1.31998,  1.32064,  1.32129,  1.32191,  1.32252,  1.32315,  1.32379,  1.32442,  1.32505,  1.32567,  1.32629,  1.32691,  1.32752,  1.32812,  1.32873,  1.32933,  1.32993,  1.33051,  1.33107,  1.33162,  1.33217,  1.33271,  1.33326,  1.33382,  1.33438,  1.33490,  1.33539,  1.33587,  1.33635,  1.33682,  1.33730,  1.33777,  1.33823,  1.33868,  1.33912,  1.33955,  1.33997,  1.34040,  1.34083,  1.34124,  1.34165,  1.34207,  1.34248,  1.34290,  1.34330,  1.34367,  1.34405,  1.34445,  1.34484,  1.34522,  1.34559,  1.34596,  1.34632,  1.34667,  1.34700,  1.34730,  1.34760,  1.34790,  1.34820,  1.34848,  1.34875,  1.34901,  1.34928,  1.34956,  1.34986,  1.35015,  1.35041,  1.35067,  1.35095,  1.35121,  1.35145,  1.35171,  1.35198,  1.35223,  1.35247,  1.35271,  1.35295,  1.35319,  1.35342,  1.35366,  1.35389,  1.35413,  1.35437,  1.35460,  1.35484,  1.35508,  1.35532,  1.35555,  1.35579,  1.35601,  1.35625,  1.35650,  1.35677,  1.35704,  1.35731,  1.35757,  1.35784,  1.35811,  1.35839,  1.35868,  1.35899,  1.35929,  1.35960,  1.35990,  1.36018,  1.36046,  1.36075,  1.36104,  1.36133,  1.36163,  1.36193,  1.36225,  1.36257,  1.36289,  1.36321,  1.36351,  1.36381,  1.36410,  1.36438,  1.36462,  1.36485,  1.36506,  1.36526,  1.36542,  1.36554,  1.36561,  1.36568,  1.36575,  1.36582,  1.36587,  1.36589,  1.36592,  1.36597,  1.36602,  1.36604,  1.36602,  1.36598,  1.36594,  1.36590,  1.36584,  1.36574,  1.36563,  1.36551,  1.36540,  1.36527,  1.36514,  1.36501,  1.36489,  1.36480,  1.36474,  1.36472,  1.36471,  1.36472,  1.36474,  1.36479,  1.36487,  1.36499,  1.36515,  1.36533,  1.36553,  1.36575,  1.36600,  1.36628,  1.36658,  1.36690,  1.36724,  1.36760,  1.36797,  1.36838,  1.36882,  1.36927,  1.36975,  1.37020,  1.37066,  1.37111,  1.37156,  1.37200,  1.37245,  1.37287,  1.37329,  1.37371,  1.37412,  1.37452,  1.37494,  1.37537,  1.37584,  1.37632,  1.37683,  1.37733,  1.37784,  1.37836,  1.37888,  1.37939,  1.37987,  1.38033,  1.38078,  1.38124,  1.38170,  1.38215,  1.38262,  1.38309,  1.38359,  1.38408,  1.38457,  1.38508,  1.38558,  1.38610,  1.38664,  1.38720,  1.38778,  1.38837,  1.38897,  1.38958,  1.39021,  1.39081,  1.39142,  1.39204,  1.39267,  1.39329,  1.39392,  1.39456,  1.39518,  1.39578,  1.39633,  1.39687,  1.39739,  1.39792,  1.39847,  1.39902,  1.39955,  1.40004,  1.40053,  1.40100,  1.40146,  1.40191,  1.40236,  1.40279,  1.40323,  1.40367,  1.40410,  1.40453,  1.40495,  1.40536,  1.40577,  1.40616,  1.40655,  1.40691,  1.40727,  1.40762,  1.40798,  1.40833,  1.40866,  1.40898,  1.40929,  1.40959,  1.40989,  1.41016,  1.41042,  1.41068,  1.41094,  1.41117,  1.41137,  1.41155,  1.41174,  1.41192,  1.41211,  1.41231,  1.41250,  1.41268,  1.41287,  1.41303,  1.41317,  1.41331,  1.41344,  1.41358,  1.41373,  1.41386,  1.41398,  1.41409,  1.41417,  1.41423,  1.41430,  1.41438,  1.41447,  1.41454,  1.41461,  1.41468,  1.41476,  1.41482,  1.41486,  1.41489,  1.41494,  1.41498,  1.41501,  1.41504,  1.41507,  1.41508,  1.41512,  1.41514,  1.41515,  1.41516,  1.41516,  1.41517,  1.41518,  1.41518,  1.41519,  1.41520,  1.41522,  1.41524,  1.41526,  1.41528,  1.41530,  1.41531,  1.41532,  1.41532,  1.41531,  1.41531,  1.41531,  1.41533,  1.41535,  1.41538,  1.41541,  1.41546,  1.41550,  1.41555,  1.41560,  1.41565,  1.41568,  1.41572,  1.41576,  1.41580,  1.41584,  1.41590,  1.41596,  1.41602,  1.41605,  1.41608,  1.41611,  1.41614,  1.41618,  1.41623,  1.41627,  1.41629,  1.41631,  1.41633,  1.41634,  1.41636,  1.41638,  1.41639,  1.41640,  1.41640,  1.41641,  1.41641,  1.41643,  1.41645,  1.41648,  1.41655,  1.41654,  1.41635,  1.41616,  1.41618,  1.41626,  1.41614,  1.41589,  1.41583,  1.41600,  1.41603,  1.41589,  1.41590,  1.41592,  1.41596,  1.41616,  1.41630,  1.41613,  1.41587,  1.41588,  1.41599,  1.41583,  1.41566,  1.41572,  1.41582,  1.41577,  1.41541,  1.41489,  1.41471,  1.41475,  1.41474,  1.41489,  1.41510,  1.41501,  1.41481,  1.41467,  1.41461,  1.41475,  1.41496,  1.41504,  1.41495,  1.41482,  1.41501,  1.41533,  1.41524,  1.41500,  1.41482,  1.41462,  1.41462,  1.41470,  1.41454,  1.41429,  1.41415,  1.41402,  1.41385,  1.41370,  1.41365,  1.41355,  1.41348,  1.41351,  1.41343,  1.41328,  1.41321,  1.41314,  1.41303,  1.41281,  1.41254,  1.41237,  1.41220,  1.41182,  1.41147,  1.41131,  1.41118,  1.41101,  1.41087,  1.41070,  1.41030,  1.40978,  1.40948,  1.40925,  1.40891,  1.40888,  1.40905,  1.40894,  1.40882,  1.40876,  1.40847,  1.40808,  1.40770,  1.40733,  1.40705,  1.40682,  1.40649,  1.40624,  1.40626,  1.40626,  1.40608,  1.40577,  1.40533,  1.40495,  1.40470,  1.40445,  1.40432,  1.40436,  1.40443,  1.40435,  1.40402,  1.40355,  1.40320,  1.40296,  1.40280,  1.40276,  1.40275,  1.40263,  1.40274,  1.40310,  1.40310,  1.40265,  1.40217,  1.40181,  1.40161,  1.40158,  1.40161,  1.40155,  1.40157,  1.40164,  1.40137,  1.40096,  1.40090,  1.40089,  1.40085,  1.40102,  1.40107,  1.40086,  1.40070,  1.40068,  1.40070,  1.40059,  1.40042,  1.40053,  1.40079,  1.40080,  1.40062,  1.40050,  1.40045,  1.40042,  1.40046,  1.40057,  1.40074,  1.40088,  1.40085,  1.40091,  1.40098,  1.40072,  1.40067,  1.40096,  1.40101,  1.40095,  1.40101,  1.40100,  1.40096,  1.40106,  1.40109,  1.40095,  1.40102,  1.40133,  1.40160,  1.40150,  1.40102,  1.40085,  1.40115,  1.40140,  1.40145,  1.40141,  1.40141,  1.40157,  1.40177,  1.40181,  1.40178,  1.40184,  1.40185,  1.40182,  1.40187,  1.40195,  1.40191,  1.40186,  1.40194,  1.40208,  1.40225,  1.40242,  1.40256,  1.40261,  1.40233,  1.40208,  1.40227,  1.40242,  1.40241,  1.40251,  1.40243,  1.40218,  1.40208,  1.40217,  1.40227,  1.40212,  1.40185,  1.40167,  1.40138,  1.40105,  1.40089,  1.40084,  1.40072,  1.40044,  1.40014,  1.39997,  1.39989,  1.39973,  1.39939,  1.39894,  1.39850,  1.39808,  1.39788,  1.39781,  1.39766,  1.39741,  1.39698,  1.39641,  1.39601,  1.39582,  1.39553,  1.39514,  1.39478,  1.39439,  1.39401,  1.39367,  1.39334,  1.39303,  1.39268,  1.39227,  1.39174,  1.39108,  1.39056,  1.39021,  1.38986,  1.38953,  1.38925,  1.38885,  1.38835,  1.38787,  1.38737,  1.38684,  1.38630,  1.38570,  1.38501,  1.38453,  1.38417,  1.38358,  1.38286,  1.38219,  1.38160,  1.38109,  1.38055,  1.37981,  1.37906,  1.37860,  1.37820,  1.37753,  1.37675,  1.37614,  1.37565,  1.37513,  1.37463,  1.37415,  1.37350,  1.37270,  1.37191,  1.37119,  1.37059,  1.36998,  1.36928,  1.36872,  1.36817,  1.36742,  1.36673,  1.36607,  1.36524,  1.36446,  1.36388,  1.36330,  1.36262,  1.36183,  1.36104,  1.36044,  1.35990,  1.35919,  1.35834,  1.35749,  1.35675,  1.35611,  1.35534,  1.35454,  1.35394,  1.35336,  1.35260,  1.35165,  1.35078,  1.35013,  1.34957,  1.34892,  1.34823,  1.34748,  1.34655,  1.34559,  1.34485,  1.34422,  1.34348,  1.34277,  1.34212,  1.34136,  1.34057,  1.33984,  1.33908,  1.33831,  1.33762,  1.33695,  1.33625,  1.33557,  1.33482,  1.33400,  1.33330,  1.33262,  1.33187,  1.33123,  1.33074,  1.33022,  1.32953,  1.32867,  1.32797,  1.32756,  1.32716,  1.32645,  1.32567,  1.32540,  1.32538,  1.32485,  1.32415,  1.32367,  1.32315,  1.32273,  1.32245,  1.32200,  1.32156,  1.32131,  1.32102,  1.32077,  1.32057,  1.32036,  1.32026,  1.32017,  1.31986,  1.31947,  1.31929,  1.31933,  1.31938,  1.31941,  1.31958,  1.31958,  1.31925,  1.31915,  1.31941,  1.31970,  1.32001,  1.32044,  1.32080,  1.32100,  1.32126,  1.32157,  1.32188,  1.32228,  1.32275,  1.32334,  1.32399,  1.32462,  1.32529,  1.32600,  1.32670,  1.32743,  1.32803,  1.32845,  1.32914,  1.33015,  1.33112,  1.33187,  1.33282,  1.33409,  1.33512,  1.33604,  1.33740,  1.33884,  1.33998,  1.34113,  1.34244,  1.34383,  1.34540,  1.34715,  1.34899,  1.35086,  1.35265,  1.35423,  1.35582,  1.35766,  1.35959,  1.36144,  1.36337,  1.36552,  1.36788,  1.37041,  1.37318,  1.37590,  1.37810,  1.38006,  1.38238,  1.38497,  1.38765,  1.39031,  1.39292,  1.39586,  1.39866,  1.40092,  1.40349,  1.40658,  1.40966,  1.41287,  1.41622,  1.41922,  1.42211,  1.42534,  1.42907,  1.43290,  1.43615,  1.43916,  1.44253,  1.44589,  1.44892,  1.45197,  1.45523,  1.45863,  1.46199,  1.46519,  1.46835,  1.47144,  1.47425,  1.47675,  1.47901,  1.48154,  1.48441,  1.48693,  1.48916,  1.49138,  1.49344,  1.49537,  1.49710,  1.49867,  1.50042,  1.50212,  1.50358,  1.50487,  1.50593,  1.50668,  1.50732,  1.50813,  1.50942,  1.51077,  1.51121,  1.51118,  1.51150,  1.51191,  1.51206,  1.51204,  1.51199,  1.51198,  1.51168,  1.51122,  1.51102,  1.51061,  1.50989,  1.50933,  1.50870,  1.50757,  1.50642,  1.50561,  1.50456,  1.50316,  1.50165,  1.49975,  1.49760,  1.49564,  1.49393,  1.49233,  1.49051,  1.48835,  1.48614,  1.48397,  1.48177,  1.47950,  1.47710,  1.47461,  1.47215,  1.46979,  1.46740,  1.46494,  1.46274,  1.46064,  1.45837,  1.45625,  1.45440,  1.45247,  1.44998,  1.44708,  1.44491,  1.44334,  1.44119,  1.43894,  1.43694,  1.43462,  1.43228,  1.43029,  1.42841,  1.42641,  1.42455,  1.42309,  1.42137,  1.41904,  1.41669,  1.41451,  1.41244,  1.41050,  1.40839,  1.40631,  1.40470,  1.40315,  1.40127,  1.39947,  1.39778,  1.39592,  1.39407,  1.39244,  1.39099,  1.38955,  1.38793,  1.38622,  1.38467,  1.38317,  1.38158,  1.38004,  1.37869,  1.37731,  1.37582,  1.37433,  1.37287,  1.37148,  1.36997,  1.36824,  1.36652,  1.36501,  1.36362,  1.36217,  1.36062,  1.35919,  1.35796,  1.35665,  1.35510,  1.35366,  1.35237,  1.35079,  1.34893,  1.34717,  1.34566,  1.34431,  1.34291,  1.34135,  1.33969,  1.33788,  1.33618,  1.33504,  1.33423,  1.33309,  1.33113,  1.32869,  1.32664,  1.32495,  1.32320,  1.32176,  1.32058,  1.31875,  1.31636,  1.31430,  1.31246,  1.31037,  1.30829,  1.30611,  1.30354,  1.30109,  1.29925,  1.29774,  1.29618,  1.29474,  1.29330,  1.29163,  1.28984,  1.28795,  1.28604,  1.28425,  1.28258,  1.28130,  1.28037,  1.27926,  1.27785,  1.27576,  1.27286,  1.27032,  1.26881,  1.26796,  1.26796,  1.26838,  1.26816,  1.26707,  1.26544,  1.26357,  1.26147,  1.25907,  1.25654,  1.25399,  1.25191,  1.25062,  1.24941,  1.24790,  1.24650,  1.24525,  1.24424,  1.24344,  1.24252,  1.24174,  1.24109,  1.24014,  1.23922,  1.23872,  1.23819,  1.23720,  1.23578,  1.23426,  1.23295,  1.23158,  1.22983,  1.22779,  1.22565,  1.22345,  1.22087,  1.21765,  1.21453,  1.21171,  1.20835,  1.20440,  1.20031,  1.19584,  1.19098,  1.18596,  1.18062,  1.17497,  1.16918,  1.16320,  1.15727,  1.15181,  1.14628,  1.14040,  1.13531,  1.13095,  1.12633,  1.12103,  1.11548,  1.11074,  1.10664,  1.10255,  1.09931,  1.09715,  1.09540,  1.09387,  1.09272,  1.09207,  1.09214,  1.09293,  1.09429,  1.09616,  1.09845,  1.10113,  1.10415,  1.10751,  1.11124,  1.11517,  1.11908,  1.12290,  1.12677,  1.13093,  1.13562,  1.14073,  1.14572,  1.15019,  1.15413,  1.15809,  1.16248,  1.16742,  1.17289,  1.17841,  1.18375,  1.18914,  1.19498,  1.20168,  1.20954,  1.21859,  1.22876,  1.23963,  1.25046,  1.26083,  1.27114,  1.28221,  1.29460,  1.30837,  1.32283,  1.33674,  1.34981,  1.36201,  1.37292,  1.38273,  1.39235,  1.40212,  1.41204,  1.42216,  1.43148,  1.43860,  1.44384,  1.44909,  1.45499,  1.46058,  1.46597,  1.47000,  1.47140,  1.47262,  1.47646,  1.48178,  1.48624,  1.49037,  1.49479,  1.49835,  1.50248,  1.50894,  1.51541,  1.51956,  1.52349,  1.52998,  1.53877,  1.54849,  1.55797,  1.56412,  1.56530,  1.56471,  1.56576,  1.56768,  1.56869,  1.56919,  1.56911,  1.56809,  1.56793,  1.56902,  1.57122,  1.57679,  1.58652,  1.59768,  1.60867,  1.62071,  1.63483,  1.65119,  1.67012,  1.69084,  1.71228,  1.73470,  1.75828,  1.78190,  1.80509,  1.82821,  1.85219,  1.87779,  1.90396,  1.92934,  1.95455,  1.97985,  2.00349,  2.02393,  2.04134,  2.05611,  2.06928,  2.08203,  2.09460,  2.10560,  2.11455,  2.12181,  2.12727,  2.13028,  2.13120,  2.13033,  2.12729,  2.12143,  2.11357,  2.10511,  2.09676,  2.08722,  2.07632,  2.06596,  2.05947,  2.05792,  2.06125,  2.06645,  2.06875,  2.06812,  2.06654,  2.06235,  2.05653,  2.05218,  2.04818,  2.04387,  2.03874,  2.03260,  2.02640,  2.02070,  2.01264,  2.00187,  1.99248,  1.98561,  1.97784,  1.96964,  1.96168,  1.95237,  1.94303,  1.93499,  1.92740,  1.91972,  1.91159,  1.90386,  1.89810,  1.89327,  1.88769,  1.88265,  1.87949,  1.87833,  1.87872,  1.88066,  1.88451,  1.89059,  1.89734,  1.90415,  1.91333,  1.92573,  1.93888,  1.95135,  1.96301,  1.97357,  1.98414,  1.99574,  2.00656,  2.01486,  2.02147,  2.02658,  2.03068,  2.03475,  2.03686,  2.03509,  2.03014,  2.02410,  2.01966,  2.01791,  2.01731,  2.01656,  2.01498,  2.01241,  2.00861,  2.00361,  1.99740,  1.99027,  1.98265,  1.97496,  1.96739,  1.96041,  1.95419,  1.94836,  1.94286,  1.93832,  1.93465,  1.93129,  1.92791,  1.92449,  1.92086,  1.91708,  
1.757,    1.741,    1.726,    1.701,    1.681,    1.663,    1.643,    1.613,    1.596,    1.551,    
1.512,    1.512,    1.542,    1.621,    1.741,    1.869,    1.939,    1.946,    1.926,    1.892,    
1.842,    1.823,    1.804,    1.782,    1.781,    1.848,    1.881,    1.918,    1.939,    1.930  ;
 
 idx_rfr_H2SO4_220K_72_NNM98_img = 
1.07e-8, 1.07e-8, 1.07e-8, 1.07e-8,
0.00E+00,  0.00E+00,  0.00E+00,  0.00E+00,  2.07E-08,  2.79E-08,  3.58E-08,  4.80E-08,  6.83E-08,  7.84E-08,  
8.20E-08,  8.39E-08,  8.46E-08,  8.79E-08,  9.98E-08,  1.24E-07,  1.58E-07,  1.83E-07,  2.02E-07,  2.33E-07,  
2.84E-07,  3.62E-07,  6.05E-07,  1.03E-06,  1.41E-06,  1.53E-06,  1.52E-06,  1.48E-06,  1.50E-06,  1.60E-06,  
1.84E-06,  2.46E-06,  4.05E-06,  4.95E-06,  5.63E-06,  6.94E-06,  7.75E-06,  8.93E-06,  1.05E-05,  1.27E-05,  
1.59E-05,  1.98E-05,  2.59E-05,  3.89E-05,  6.16E-05,  8.78E-05,  1.02E-04,  1.10E-04,  1.17E-04,  1.25E-04,  
1.38E-04,  1.55E-04,  1.76E-04,  2.02E-04,  2.34E-04,  2.72E-04,  3.14E-04,  3.61E-04,  4.24E-04,  4.86E-04,  
5.37E-04,  5.95E-04,  7.96E-04,  1.11E-03,  1.24E-03,  1.26E-03,  1.30E-03,  1.35E-03,
 0.00198,  0.00207,  0.00126,  0.00027,  0.00143,  0.00168,  0.00027,  0.00003,  0.00054,  0.00036,  0.00087,  0.00135,  0.00027,  0.00034,  0.00075,  0.00132,  0.00167,  0.00148,  0.00110,  0.00082,  0.00008,  0.00049,  0.00174,  0.00240,  0.00177,  0.00161,  0.00153,  0.00111,  0.00143,  0.00114,  0.00071,  0.00092,  0.00207,  0.00204,  0.00038,  0.00029,  0.00097,  0.00118,  0.00118,  0.00127,  0.00170,  0.00112,  0.00080,  0.00037,  0.00008,  0.00001,  0.00094,  0.00218,  0.00131,  0.00099,  0.00037,  0.00124,  0.00107,  0.00053,  0.00096,  0.00022,  0.00076,  0.00005,  0.00033,  0.00016,  0.00015,  0.00017,  0.00101,  0.00094,  0.00084,  0.00183,  0.00148,  0.00084,  0.00082,  0.00107,  0.00167,  0.00074,  0.00023,  0.00116,  0.00098,  0.00006,  0.00112,  0.00109,  0.00008,  0.00008,  0.00003,  0.00075,  0.00058,  0.00052,  0.00115,  0.00055,  0.00114,  0.00012,  0.00098,  0.00124,  0.00085,  0.00120,  0.00153,  0.00093,  0.00021,  0.00017,  0.00013,  0.00055,  0.00006,  0.00116,  0.00113,  0.00012,  0.00049,  0.00002,  0.00095,  0.00022,  0.00044,  0.00106,  0.00001,  0.00137,  0.00122,  0.00129,  0.00128,  0.00070,  0.00075,  0.00095,  0.00082,  0.00010,  0.00052,  0.00035,  0.00077,  0.00062,  0.00037,  0.00050,  0.00124,  0.00062,  0.00048,  0.00023,  0.00004,  0.00027,  0.00099,  0.00101,  0.00003,  0.00074,  0.00078,  0.00071,  0.00167,  0.00130,  0.00065,  0.00093,  0.00101,  0.00086,  0.00075,  0.00038,  0.00034,  0.00018,  0.00038,  0.00169,  0.00238,  0.00267,  0.00179,  0.00122,  0.00135,  0.00155,  0.00074,  0.00037,  0.00010,  0.00022,  0.00242,  0.00241,  0.00050,  0.00095,  0.00156,  0.00092,  0.00116,  0.00231,  0.00192,  0.00167,  0.00139,  0.00000,  0.00030,  0.00049,  0.00094,  0.00164,  0.00303,  0.00397,  0.00305,  0.00159,  0.00116,  0.00108,  0.00074,  0.00100,  0.00189,  0.00108,  0.00038,  0.00050,  0.00104,  0.00153,  0.00104,  0.00192,  0.00263,  0.00165,  0.00073,  0.00177,  0.00400,  0.00329,  0.00146,  0.00160,  0.00158,  0.00147,  0.00056,  0.00041,  0.00150,  0.00301,  0.00365,  0.00202,  0.00215,  0.00229,  0.00164,  0.00288,  0.00373,  0.00383,  0.00287,  0.00180,  0.00193,  0.00171,  0.00204,  0.00240,  0.00203,  0.00127,  0.00060,  0.00103,  0.00195,  0.00254,  0.00215,  0.00138,  0.00165,  0.00238,  0.00261,  0.00240,  0.00246,  0.00222,  0.00213,  0.00339,  0.00349,  0.00295,  0.00238,  0.00222,  0.00293,  0.00221,  0.00124,  0.00172,  0.00223,  0.00196,  0.00174,  0.00191,  0.00208,  0.00141,  0.00123,  0.00241,  0.00220,  0.00121,  0.00153,  0.00180,  0.00163,  0.00138,  0.00154,  0.00203,  0.00208,  0.00216,  0.00153,  0.00179,  0.00292,  0.00213,  0.00084,  0.00090,  0.00183,  0.00238,  0.00254,  0.00233,  0.00197,  0.00151,  0.00137,  0.00261,  0.00296,  0.00256,  0.00343,  0.00383,  0.00273,  0.00240,  0.00284,  0.00228,  0.00160,  0.00185,  0.00201,  0.00210,  0.00263,  0.00297,  0.00301,  0.00251,  0.00241,  0.00314,  0.00322,  0.00324,  0.00308,  0.00260,  0.00242,  0.00192,  0.00174,  0.00246,  0.00265,  0.00212,  0.00191,  0.00194,  0.00208,  0.00288,  0.00305,  0.00240,  0.00232,  0.00205,  0.00171,  0.00194,  0.00197,  0.00205,  0.00130,  0.00165,  0.00295,  0.00266,  0.00246,  0.00238,  0.00282,  0.00366,  0.00337,  0.00234,  0.00215,  0.00196,  0.00134,  0.00181,  0.00243,  0.00242,  0.00244,  0.00288,  0.00270,  0.00229,  0.00185,  0.00167,  0.00179,  0.00168,  0.00153,  0.00126,  0.00189,  0.00246,  0.00213,  0.00262,  0.00315,  0.00294,  0.00308,  0.00355,  0.00370,  0.00424,  0.00414,  0.00318,  0.00268,  0.00238,  0.00301,  0.00332,  0.00347,  0.00348,  0.00230,  0.00218,  0.00223,  0.00228,  0.00286,  0.00189,  0.00189,  0.00306,  0.00318,  0.00363,  0.00340,  0.00266,  0.00284,  0.00311,  0.00297,  0.00317,  0.00334,  0.00321,  0.00359,  0.00377,  0.00322,  0.00309,  0.00301,  0.00291,  0.00335,  0.00260,  0.00139,  0.00125,  0.00221,  0.00318,  0.00252,  0.00191,  0.00267,  0.00315,  0.00216,  0.00184,  0.00310,  0.00284,  0.00211,  0.00271,  0.00302,  0.00269,  0.00277,  0.00255,  0.00142,  0.00127,  0.00204,  0.00265,  0.00293,  0.00292,  0.00320,  0.00304,  0.00227,  0.00284,  0.00344,  0.00304,  0.00243,  0.00185,  0.00193,  0.00248,  0.00329,  0.00351,  0.00303,  0.00267,  0.00263,  0.00269,  0.00267,  0.00259,  0.00260,  0.00248,  0.00281,  0.00331,  0.00324,  0.00325,  0.00316,  0.00299,  0.00275,  0.00292,  0.00344,  0.00308,  0.00269,  0.00304,  0.00306,  0.00306,  0.00299,  0.00275,  0.00292,  0.00283,  0.00230,  0.00208,  0.00205,  0.00203,  0.00260,  0.00299,  0.00282,  0.00285,  0.00303,  0.00273,  0.00267,  0.00321,  0.00317,  0.00292,  0.00259,  0.00226,  0.00184,  0.00159,  0.00223,  0.00228,  0.00199,  0.00229,  0.00220,  0.00183,  0.00192,  0.00238,  0.00290,  0.00264,  0.00171,  0.00162,  0.00235,  0.00241,  0.00193,  0.00172,  0.00199,  0.00215,  0.00202,  0.00164,  0.00105,  0.00096,  0.00180,  0.00223,  0.00175,  0.00223,  0.00236,  0.00183,  0.00227,  0.00267,  0.00236,  0.00179,  0.00136,  0.00142,  0.00157,  0.00190,  0.00218,  0.00189,  0.00166,  0.00190,  0.00195,  0.00157,  0.00164,  0.00226,  0.00230,  0.00161,  0.00129,  0.00189,  0.00208,  0.00157,  0.00148,  0.00182,  0.00199,  0.00188,  0.00145,  0.00133,  0.00099,  0.00070,  0.00118,  0.00087,  0.00018,  0.00053,  0.00072,  0.00017,  0.00038,  0.00066,  0.00030,  0.00022,  0.00006,  0.00046,  0.00075,  0.00076,  0.00066,  0.00108,  0.00104,  0.00074,  0.00097,  0.00126,  0.00173,  0.00189,  0.00236,  0.00315,  0.00357,  0.00372,  0.00388,  0.00432,  0.00459,  0.00505,  0.00523,  0.00530,  0.00584,  0.00671,  0.00740,  0.00762,  0.00796,  0.00852,  0.00935,  0.00971,  0.01025,  0.01129,  0.01172,  0.01210,  0.01278,  0.01356,  0.01428,  0.01515,  0.01559,  0.01609,  0.01737,  0.01812,  0.01912,  0.02026,  0.02057,  0.02117,  0.02206,  0.02328,  0.02459,  0.02548,  0.02576,  0.02595,  0.02765,  0.02920,  0.02994,  0.03106,  0.03216,  0.03314,  0.03343,  0.03351,  0.03460,  0.03630,  0.03764,  0.03865,  0.03984,  0.04126,  0.04216,  0.04215,  0.04300,  0.04392,  0.04453,  0.04545,  0.04614,  0.04681,  0.04743,  0.04865,  0.05042,  0.05294,  0.05414,  0.05398,  0.05490,  0.05601,  0.05657,  0.05710,  0.05796,  0.05864,  0.06026,  0.06167,  0.06205,  0.06346,  0.06418,  0.06521,  0.06678,  0.06668,  0.06721,  0.06848,  0.07023,  0.07156,  0.07171,  0.07161,  0.07225,  0.07386,  0.07512,  0.07604,  0.07666,  0.07795,  0.07844,  0.07868,  0.07983,  0.08028,  0.08084,  0.08204,  0.08394,  0.08508,  0.08494,  0.08591,  0.08724,  0.08859,  0.08966,  0.08918,  0.09012,  0.09155,  0.09137,  0.09143,  0.09277,  0.09390,  0.09449,  0.09558,  0.09642,  0.09679,  0.09643,  0.09689,  0.09848,  0.09910,  0.10010,  0.10124,  0.10051,  0.10094,  0.10263,  0.10279,  0.10317,  0.10359,  0.10420,  0.10592,  0.10649,  0.10617,  0.10670,  0.10701,  0.10654,  0.10703,  0.10757,  0.10766,  0.10855,  0.11014,  0.11150,  0.11113,  0.11085,  0.11248,  0.11362,  0.11347,  0.11288,  0.11299,  0.11364,  0.11412,  0.11461,  0.11462,  0.11429,  0.11417,  0.11388,  0.11368,  0.11527,  0.11657,  0.11673,  0.11700,  0.11802,  0.11864,  0.11883,  0.11917,  0.11835,  0.11871,  0.11891,  0.11898,  0.11990,  0.11910,  0.11843,  0.11939,  0.12086,  0.12027,  0.11870,  0.11920,  0.11999,  0.12150,  0.12262,  0.12180,  0.12112,  0.12133,  0.12221,  0.12276,  0.12245,  0.12248,  0.12281,  0.12366,  0.12488,  0.12345,  0.12236,  0.12413,  0.12471,  0.12372,  0.12439,  0.12558,  0.12530,  0.12497,  0.12537,  0.12497,  0.12511,  0.12609,  0.12667,  0.12687,  0.12670,  0.12674,  0.12558,  0.12574,  0.12648,  0.12688,  0.12827,  0.12864,  0.12892,  0.12911,  0.12906,  0.13031,  0.13155,  0.13111,  0.13149,  0.13193,  0.13100,  0.13070,  0.13142,  0.13237,  0.13315,  0.13395,  0.13331,  0.13300,  0.13368,  0.13328,  0.13398,  0.13446,  0.13499,  0.13545,  0.13464,  0.13532,  0.13593,  0.13549,  0.13431,  0.13317,  0.13397,  0.13586,  0.13714,  0.13712,  0.13619,  0.13592,  0.13686,  0.13796,  0.13849,  0.13851,  0.13877,  0.13912,  0.13941,  0.13966,  0.13989,  0.14071,  0.14074,  0.14082,  0.14090,  0.14042,  0.14071,  0.13983,  0.14004,  0.14165,  0.14208,  0.14197,  0.14180,  0.14246,  0.14386,  0.14453,  0.14324,  0.14245,  0.14388,  0.14505,  0.14542,  0.14520,  0.14404,  0.14489,  0.14711,  0.14777,  0.14832,  0.14859,  0.14727,  0.14603,  0.14656,  0.14725,  0.14798,  0.14839,  0.14811,  0.14904,  0.15016,  0.15008,  0.14938,  0.14999,  0.15036,  0.15045,  0.15161,  0.15213,  0.15230,  0.15208,  0.15208,  0.15232,  0.15209,  0.15229,  0.15353,  0.15411,  0.15441,  0.15597,  0.15608,  0.15525,  0.15594,  0.15697,  0.15732,  0.15648,  0.15556,  0.15635,  0.15715,  0.15709,  0.15660,  0.15710,  0.15907,  0.15946,  0.15933,  0.16012,  0.16043,  0.16086,  0.16169,  0.16192,  0.16182,  0.16236,  0.16285,  0.16333,  0.16385,  0.16368,  0.16341,  0.16370,  0.16376,  0.16353,  0.16426,  0.16445,  0.16435,  0.16471,  0.16493,  0.16552,  0.16580,  0.16495,  0.16483,  0.16608,  0.16591,  0.16517,  0.16491,  0.16444,  0.16420,  0.16413,  0.16438,  0.16557,  0.16618,  0.16519,  0.16431,  0.16464,  0.16569,  0.16641,  0.16665,  0.16670,  0.16703,  0.16635,  0.16570,  0.16574,  0.16574,  0.16616,  0.16600,  0.16577,  0.16624,  0.16737,  0.16885,  0.16960,  0.16969,  0.17081,  0.17263,  0.17216,  0.17113,  0.17257,  0.17349,  0.17304,  0.17267,  0.17345,  0.17410,  0.17314,  0.17324,  0.17400,  0.17406,  0.17331,  0.17320,  0.17423,  0.17359,  0.17235,  0.17173,  0.17172,  0.17243,  0.17256,  0.17252,  0.17331,  0.17389,  0.17283,  0.17245,  0.17301,  0.17285,  0.17299,  0.17290,  0.17316,  0.17426,  0.17477,  0.17491,  0.17472,  0.17483,  0.17537,  0.17541,  0.17529,  0.17473,  0.17541,  0.17607,  0.17512,  0.17546,  0.17574,  0.17517,  0.17546,  0.17511,  0.17407,  0.17431,  0.17374,  0.17270,  0.17317,  0.17393,  0.17395,  0.17283,  0.17294,  0.17331,  0.17211,  0.17147,  0.17148,  0.17093,  0.17128,  0.17162,  0.17043,  0.17018,  0.16992,  0.16979,  0.17066,  0.17101,  0.17056,  0.17008,  0.16966,  0.16968,  0.16943,  0.16820,  0.16780,  0.16748,  0.16734,  0.16768,  0.16750,  0.16699,  0.16693,  0.16647,  0.16558,  0.16547,  0.16538,  0.16487,  0.16398,  0.16402,  0.16443,  0.16417,  0.16312,  0.16245,  0.16285,  0.16299,  0.16315,  0.16272,  0.16206,  0.16205,  0.16162,  0.16095,  0.15996,  0.15950,  0.15976,  0.15924,  0.15839,  0.15813,  0.15863,  0.15797,  0.15692,  0.15695,  0.15672,  0.15684,  0.15695,  0.15670,  0.15624,  0.15619,  0.15700,  0.15622,  0.15542,  0.15568,  0.15554,  0.15547,  0.15492,  0.15468,  0.15493,  0.15452,  0.15375,  0.15337,  0.15270,  0.15232,  0.15299,  0.15360,  0.15362,  0.15320,  0.15255,  0.15196,  0.15225,  0.15190,  0.15106,  0.15121,  0.15207,  0.15278,  0.15258,  0.15194,  0.15105,  0.15104,  0.15135,  0.15075,  0.15028,  0.15007,  0.14992,  0.15027,  0.15033,  0.15025,  0.14997,  0.15006,  0.15056,  0.15067,  0.15072,  0.15006,  0.14930,  0.14907,  0.15006,  0.15048,  0.14945,  0.14917,  0.14919,  0.14901,  0.14924,  0.14922,  0.14867,  0.14847,  0.14842,  0.14832,  0.14885,  0.14949,  0.14897,  0.14885,  0.14899,  0.14867,  0.14841,  0.14774,  0.14773,  0.14825,  0.14828,  0.14805,  0.14770,  0.14744,  0.14728,  0.14681,  0.14685,  0.14737,  0.14719,  0.14637,  0.14610,  0.14646,  0.14661,  0.14695,  0.14716,  0.14712,  0.14677,  0.14620,  0.14625,  0.14588,  0.14551,  0.14595,  0.14600,  0.14521,  0.14442,  0.14448,  0.14480,  0.14484,  0.14494,  0.14474,  0.14400,  0.14378,  0.14372,  0.14371,  0.14426,  0.14424,  0.14368,  0.14352,  0.14374,  0.14382,  0.14395,  0.14406,  0.14421,  0.14429,  0.14372,  0.14329,  0.14264,  0.14176,  0.14120,  0.14130,  0.14136,  0.14032,  0.13949,  0.13964,  0.13998,  0.14044,  0.14103,  0.14044,  0.13941,  0.13903,  0.13902,  0.13916,  0.13890,  0.13819,  0.13770,  0.13792,  0.13764,  0.13764,  0.13795,  0.13733,  0.13700,  0.13623,  0.13524,  0.13583,  0.13644,  0.13610,  0.13572,  0.13495,  0.13396,  0.13391,  0.13431,  0.13379,  0.13326,  0.13346,  0.13350,  0.13258,  0.13193,  0.13267,  0.13287,  0.13227,  0.13181,  0.13185,  0.13198,  0.13176,  0.13155,  0.13149,  0.13209,  0.13267,  0.13272,  0.13238,  0.13238,  0.13231,  0.13215,  0.13222,  0.13184,  0.13175,  0.13152,  0.13109,  0.13022,  0.12946,  0.13031,  0.13111,  0.13133,  0.13152,  0.13158,  0.13221,  0.13162,  0.13039,  0.13109,  0.13177,  0.13161,  0.13175,  0.13188,  0.13154,  0.13073,  0.13027,  0.13066,  0.13096,  0.13108,  0.13172,  0.13204,  0.13181,  0.13213,  0.13218,  0.13220,  0.13248,  0.13208,  0.13221,  0.13291,  0.13357,  0.13391,  0.13412,  0.13402,  0.13348,  0.13362,  0.13476,  0.13564,  0.13508,  0.13481,  0.13547,  0.13610,  0.13588,  0.13547,  0.13594,  0.13590,  0.13547,  0.13610,  0.13735,  0.13722,  0.13626,  0.13679,  0.13709,  0.13613,  0.13651,  0.13705,  0.13721,  0.13802,  0.13803,  0.13773,  0.13766,  0.13756,  0.13769,  0.13793,  0.13773,  0.13748,  0.13788,  0.13846,  0.13808,  0.13769,  0.13771,  0.13765,  0.13815,  0.13853,  0.13847,  0.13804,  0.13782,  0.13728,  0.13714,  0.13757,  0.13736,  0.13706,  0.13678,  0.13680,  0.13657,  0.13617,  0.13622,  0.13619,  0.13576,  0.13546,  0.13516,  0.13465,  0.13417,  0.13398,  0.13424,  0.13391,  0.13301,  0.13292,  0.13322,  0.13292,  0.13263,  0.13268,  0.13265,  0.13164,  0.13075,  0.13065,  0.13042,  0.13021,  0.13044,  0.13090,  0.13008,  0.12917,  0.12937,  0.12930,  0.12925,  0.12940,  0.12926,  0.12879,  0.12793,  0.12758,  0.12791,  0.12792,  0.12775,  0.12771,  0.12736,  0.12696,  0.12695,  0.12676,  0.12580,  0.12493,  0.12470,  0.12528,  0.12555,  0.12496,  0.12442,  0.12397,  0.12459,  0.12487,  0.12397,  0.12356,  0.12396,  0.12390,  0.12280,  0.12225,  0.12292,  0.12324,  0.12269,  0.12268,  0.12254,  0.12212,  0.12231,  0.12222,  0.12248,  0.12278,  0.12243,  0.12242,  0.12256,  0.12272,  0.12237,  0.12194,  0.12194,  0.12119,  0.12095,  0.12195,  0.12251,  0.12255,  0.12247,  0.12281,  0.12293,  0.12251,  0.12252,  0.12215,  0.12121,  0.12169,  0.12342,  0.12413,  0.12421,  0.12404,  0.12377,  0.12398,  0.12398,  0.12349,  0.12352,  0.12448,  0.12521,  0.12570,  0.12631,  0.12636,  0.12644,  0.12666,  0.12652,  0.12646,  0.12757,  0.12830,  0.12785,  0.12780,  0.12824,  0.12909,  0.12926,  0.12948,  0.13062,  0.13159,  0.13222,  0.13281,  0.13283,  0.13276,  0.13364,  0.13492,  0.13597,  0.13697,  0.13722,  0.13652,  0.13628,  0.13674,  0.13769,  0.13797,  0.13926,  0.14166,  0.14097,  0.13997,  0.14133,  0.14309,  0.14390,  0.14473,  0.14565,  0.14604,  0.14702,  0.14817,  0.14947,  0.15020,  0.15038,  0.15062,  0.15177,  0.15321,  0.15426,  0.15583,  0.15671,  0.15670,  0.15762,  0.16018,  0.16098,  0.16026,  0.16122,  0.16334,  0.16517,  0.16610,  0.16722,  0.16823,  0.16896,  0.17032,  0.17148,  0.17328,  0.17504,  0.17603,  0.17768,  0.17866,  0.17957,  0.18179,  0.18333,  0.18408,  0.18557,  0.18727,  0.18845,  0.18915,  0.19035,  0.19223,  0.19416,  0.19564,  0.19711,  0.19907,  0.20039,  0.20182,  0.20362,  0.20510,  0.20709,  0.20908,  0.21012,  0.21060,  0.21186,  0.21420,  0.21622,  0.21727,  0.21855,  0.22051,  0.22203,  0.22419,  0.22638,  0.22784,  0.23006,  0.23161,  0.23308,  0.23539,  0.23707,  0.23822,  0.23970,  0.24193,  0.24321,  0.24427,  0.24696,  0.24861,  0.24952,  0.25124,  0.25201,  0.25296,  0.25433,  0.25509,  0.25680,  0.25875,  0.25918,  0.25989,  0.26197,  0.26327,  0.26433,  0.26618,  0.26741,  0.26750,  0.26770,  0.26954,  0.27183,  0.27278,  0.27435,  0.27612,  0.27662,  0.27708,  0.27735,  0.27775,  0.27888,  0.27930,  0.27870,  0.27903,  0.27904,  0.27866,  0.27879,  0.27805,  0.27734,  0.27707,  0.27653,  0.27526,  0.27437,  0.27373,  0.27149,  0.26916,  0.26769,  0.26734,  0.26718,  0.26435,  0.26107,  0.25956,  0.25751,  0.25503,  0.25332,  0.25107,  0.24818,  0.24534,  0.24341,  0.24172,  0.23959,  0.23742,  0.23512,  0.23280,  0.23048,  0.22798,  0.22468,  0.22138,  0.21903,  0.21742,  0.21449,  0.21048,  0.20796,  0.20585,  0.20296,  0.20096,  0.19907,  0.19538,  0.19230,  0.19078,  0.18842,  0.18478,  0.18203,  0.18075,  0.17831,  0.17493,  0.17322,  0.17160,  0.16904,  0.16617,  0.16382,  0.16284,  0.16098,  0.15889,  0.15710,  0.15438,  0.15296,  0.15216,  0.15083,  0.14979,  0.14875,  0.14685,  0.14447,  0.14342,  0.14337,  0.14272,  0.14054,  0.14010,  0.14047,  0.13891,  0.13861,  0.13855,  0.13735,  0.13744,  0.13745,  0.13659,  0.13701,  0.13674,  0.13538,  0.13534,  0.13649,  0.13686,  0.13667,  0.13699,  0.13643,  0.13511,  0.13436,  0.13457,  0.13499,  0.13547,  0.13592,  0.13573,  0.13593,  0.13696,  0.13761,  0.13675,  0.13609,  0.13746,  0.13918,  0.13917,  0.13903,  0.14021,  0.14002,  0.13961,  0.14069,  0.14177,  0.14256,  0.14220,  0.14121,  0.14182,  0.14200,  0.14227,  0.14393,  0.14398,  0.14436,  0.14527,  0.14569,  0.14550,  0.14569,  0.14782,  0.14841,  0.14828,  0.14973,  0.15052,  0.15013,  0.15098,  0.15240,  0.15372,  0.15484,  0.15476,  0.15741,  0.15861,  0.15749,  0.15925,  0.16044,  0.16048,  0.16146,  0.16315,  0.16327,  0.16468,  0.16604,  0.16585,  0.16614,  0.16583,  0.16809,  0.17004,  0.16911,  0.17008,  0.17195,  0.17226,  0.17257,  0.17141,  0.17171,  0.17446,  0.17520,  0.17585,  0.17711,  0.17812,  0.17917,  0.18045,  0.18282,  0.18509,  0.18499,  0.18511,  0.18714,  0.18826,  0.18933,  0.19301,  0.19738,  0.19967,  0.20063,  0.20295,  0.20629,  0.20967,  0.21385,  0.21725,  0.22055,  0.22351,  0.22673,  0.23019,  0.23317,  0.23656,  0.23969,  0.24065,  0.24138,  0.24577,  0.25096,  0.25449,  0.25740,  0.26089,  0.26484,  0.26889,  0.27341,  0.27773,  0.28068,  0.28380,  0.28875,  0.29257,  0.29575,  0.29904,  0.30237,  0.30648,  0.30888,  0.31141,  0.31559,  0.31913,  0.32177,  0.32359,  0.32558,  0.32713,  0.32857,  0.33134,  0.33266,  0.33308,  0.33571,  0.33895,  0.34011,  0.34172,  0.34524,  0.34662,  0.34749,  0.35049,  0.35467,  0.35832,  0.36147,  0.36583,  0.37054,  0.37668,  0.38363,  0.39092,  0.39855,  0.40491,  0.41205,  0.42066,  0.42933,  0.43848,  0.44737,  0.45698,  0.46904,  0.48059,  0.49099,  0.50226,  0.51463,  0.52595,  0.53656,  0.54797,  0.55990,  0.57213,  0.58218,  0.59156,  0.60178,  0.61155,  0.62135,  0.62924,  0.63607,  0.64561,  0.65427,  0.66017,  0.66836,  0.67598,  0.68201,  0.68905,  0.69516,  0.70078,  0.70525,  0.70958,  0.71615,  0.72422,  0.73010,  0.73506,  0.74281,  0.74941,  0.75646,  0.76458,  0.76969,  0.77454,  0.78081,  0.78786,  0.79400,  0.79692,  0.79822,  0.80227,  0.80753,  0.80928,  0.80715,  0.80602,  0.80756,  0.80748,  0.80533,  0.80021,  0.79458,  0.78673,  0.77829,  0.77145,  0.76031,  0.75451,  0.75075,  0.74070,  0.73343,  0.72895,  0.71655,  0.70201,  0.70224,  0.70300,  0.69393,  0.68403,  0.67187,  0.66669,  0.66648,  0.66381,  0.66065,  0.65578,  0.65474,  0.65638,  0.65394,  0.64835,  0.64271,  0.63860,  0.63927,  0.63950,  0.63906,  0.63947,  0.64612,  0.65634,  0.65833,  0.66875,  0.68660,  0.69673,  0.70560,  0.71293,  0.72674,  0.74768,  0.76301,  0.77158,  0.77948,  0.79185,  0.79958,  0.80770,  0.81713,  0.82322,  0.82572,  0.82364,  0.82384,  0.82099,  0.81412,  0.80953,  0.79978,  0.78625,  0.77777,  0.76518,  0.74759,  0.73415,  0.71945,  0.69913,  0.68247,  0.66782,  0.65081,  0.63410,  0.61645,  0.60196,  0.58782,  0.57026,  0.55422,  0.54021,  0.52720,  0.51480,  0.50317,  0.49448,  0.48673,  0.47756,  0.47034,  0.46490,  0.46135,  0.46021,  0.45251,  0.44198,  0.43524,  0.42534,  0.41821,  0.41220,  0.40243,  0.40178,  0.39891,  0.38782,  0.38077,  0.37989,  0.37713,  0.37115,  0.36797,  0.36322,  0.36297,  0.36302,  0.35897,  0.35780,  0.35778,  0.35948,  0.35916,  0.35914,  0.36394,  0.37092,  0.37809,  0.38292,  0.38941,  0.40431,  0.41993,  0.43093,  0.44206,  0.45418,  0.46692,  0.47937,  0.49213,  0.50272,  0.51362,  0.52463,  0.52793,  0.52537,  0.52240,  0.51992,  0.51703,  0.51146,  0.50010,  0.48831,  0.47653,  0.46171,  0.44720,  0.43176,  0.41439,  0.39775,  0.38112,  0.36557,  0.35407,  0.34155,  0.32913,  0.31693,  0.30505,  0.29361,  0.28271,  0.27247,  0.26298,  0.25436,  0.24672,  0.24025,  0.23478,  0.23001,  0.22571,  0.22162,  0.21811,  0.21514,  0.21208,  0.20896,  0.20585,  0.20277,  0.19980,  0.19697,  
0.158,    0.157,    0.157,    0.16,     0.165,    0.171,    0.173,    0.183,    0.191,    0.221,    
0.299,    0.352,    0.479,    0.564,    0.594,    0.554,    0.457,    0.362,    0.299,    0.261,    
0.238,    0.235,    0.24,     0.257,    0.29,     0.329,    0.32,     0.3,      0.226,    0.2  ;

 idx_rfr_H2SO4_220K_72_NNM98_rl =
1.526, 1.512, 1.496, 1.484,
1.452,  1.438,  1.432,  1.431,  1.428,  1.427,  1.427,  1.427,  1.427,  1.427,  
1.427,  1.427,  1.427,  1.427,  1.427,  1.426,  1.426,  1.425,  1.425,  1.425,  
1.424,  1.424,  1.423,  1.423,  1.422,  1.422,  1.421,  1.421,  1.420,  1.419,  
1.418,  1.417,  1.416,  1.416,  1.415,  1.413,  1.413,  1.412,  1.411,  1.411,  
1.410,  1.410,  1.409,  1.408,  1.407,  1.406,  1.406,  1.405,  1.404,  1.403,  
1.403,  1.402,  1.400,  1.399,  1.398,  1.398,  1.397,  1.396,  1.394,  1.393,  
1.392,  1.391,  1.389,  1.388,  1.386,  1.384,  1.382,  1.380, 
 1.37992,  1.38016,  1.38033,  1.37953,  1.37904,  1.37979,  1.37991,  1.37905,  1.37862,  1.37834,  1.37815,  1.37857,  1.37862,  1.37792,  1.37744,  1.37746,  1.37782,  1.37823,  1.37834,  1.37830,  1.37767,  1.37670,  1.37649,  1.37733,  1.37784,  1.37790,  1.37789,  1.37778,  1.37768,  1.37782,  1.37746,  1.37680,  1.37702,  1.37810,  1.37811,  1.37714,  1.37666,  1.37683,  1.37682,  1.37681,  1.37711,  1.37746,  1.37743,  1.37718,  1.37672,  1.37585,  1.37536,  1.37604,  1.37682,  1.37685,  1.37622,  1.37616,  1.37638,  1.37642,  1.37623,  1.37620,  1.37604,  1.37593,  1.37562,  1.37543,  1.37513,  1.37459,  1.37456,  1.37471,  1.37449,  1.37468,  1.37531,  1.37531,  1.37485,  1.37465,  1.37511,  1.37542,  1.37476,  1.37456,  1.37499,  1.37457,  1.37428,  1.37485,  1.37487,  1.37427,  1.37371,  1.37366,  1.37367,  1.37353,  1.37352,  1.37363,  1.37370,  1.37339,  1.37303,  1.37322,  1.37333,  1.37312,  1.37362,  1.37398,  1.37380,  1.37323,  1.37288,  1.37274,  1.37234,  1.37232,  1.37288,  1.37291,  1.37246,  1.37207,  1.37211,  1.37201,  1.37173,  1.37176,  1.37150,  1.37118,  1.37151,  1.37178,  1.37195,  1.37198,  1.37160,  1.37168,  1.37184,  1.37159,  1.37117,  1.37098,  1.37093,  1.37102,  1.37081,  1.37041,  1.37064,  1.37090,  1.37083,  1.37054,  1.37017,  1.36957,  1.36967,  1.37009,  1.36983,  1.36935,  1.36932,  1.36905,  1.36922,  1.36976,  1.36962,  1.36926,  1.36930,  1.36933,  1.36931,  1.36907,  1.36875,  1.36819,  1.36741,  1.36709,  1.36769,  1.36863,  1.36916,  1.36889,  1.36858,  1.36886,  1.36891,  1.36853,  1.36773,  1.36659,  1.36674,  1.36819,  1.36820,  1.36726,  1.36731,  1.36726,  1.36664,  1.36687,  1.36745,  1.36775,  1.36796,  1.36751,  1.36651,  1.36586,  1.36532,  1.36480,  1.36503,  1.36638,  1.36776,  1.36783,  1.36723,  1.36684,  1.36636,  1.36579,  1.36609,  1.36649,  1.36602,  1.36512,  1.36476,  1.36483,  1.36456,  1.36423,  1.36490,  1.36544,  1.36445,  1.36323,  1.36409,  1.36578,  1.36585,  1.36506,  1.36491,  1.36503,  1.36455,  1.36336,  1.36232,  1.36262,  1.36394,  1.36432,  1.36384,  1.36368,  1.36315,  1.36259,  1.36316,  1.36429,  1.36490,  1.36457,  1.36402,  1.36364,  1.36339,  1.36358,  1.36402,  1.36390,  1.36307,  1.36206,  1.36176,  1.36226,  1.36275,  1.36238,  1.36163,  1.36147,  1.36179,  1.36189,  1.36191,  1.36172,  1.36115,  1.36115,  1.36193,  1.36245,  1.36226,  1.36183,  1.36203,  1.36247,  1.36192,  1.36115,  1.36119,  1.36137,  1.36114,  1.36092,  1.36110,  1.36097,  1.36020,  1.36013,  1.36076,  1.36056,  1.35994,  1.35987,  1.35992,  1.35957,  1.35915,  1.35901,  1.35915,  1.35935,  1.35907,  1.35847,  1.35885,  1.35966,  1.35918,  1.35796,  1.35742,  1.35758,  1.35796,  1.35818,  1.35820,  1.35775,  1.35683,  1.35648,  1.35689,  1.35681,  1.35676,  1.35758,  1.35798,  1.35753,  1.35749,  1.35770,  1.35722,  1.35659,  1.35628,  1.35594,  1.35574,  1.35591,  1.35626,  1.35620,  1.35570,  1.35554,  1.35582,  1.35609,  1.35632,  1.35635,  1.35625,  1.35594,  1.35526,  1.35495,  1.35527,  1.35534,  1.35498,  1.35452,  1.35405,  1.35404,  1.35456,  1.35475,  1.35461,  1.35445,  1.35409,  1.35370,  1.35357,  1.35362,  1.35311,  1.35221,  1.35220,  1.35270,  1.35265,  1.35222,  1.35191,  1.35231,  1.35313,  1.35318,  1.35280,  1.35256,  1.35197,  1.35121,  1.35111,  1.35120,  1.35105,  1.35114,  1.35146,  1.35155,  1.35126,  1.35082,  1.35049,  1.35031,  1.35001,  1.34931,  1.34875,  1.34876,  1.34861,  1.34823,  1.34833,  1.34840,  1.34814,  1.34806,  1.34811,  1.34848,  1.34917,  1.34943,  1.34899,  1.34825,  1.34782,  1.34783,  1.34812,  1.34858,  1.34852,  1.34788,  1.34735,  1.34700,  1.34711,  1.34690,  1.34594,  1.34553,  1.34572,  1.34601,  1.34638,  1.34619,  1.34566,  1.34552,  1.34539,  1.34520,  1.34517,  1.34503,  1.34496,  1.34528,  1.34540,  1.34521,  1.34500,  1.34480,  1.34504,  1.34544,  1.34488,  1.34352,  1.34274,  1.34314,  1.34356,  1.34294,  1.34240,  1.34286,  1.34290,  1.34197,  1.34173,  1.34219,  1.34183,  1.34130,  1.34145,  1.34151,  1.34150,  1.34171,  1.34130,  1.34013,  1.33934,  1.33924,  1.33935,  1.33932,  1.33942,  1.33963,  1.33919,  1.33859,  1.33880,  1.33925,  1.33915,  1.33851,  1.33762,  1.33698,  1.33699,  1.33746,  1.33768,  1.33740,  1.33701,  1.33675,  1.33656,  1.33631,  1.33604,  1.33560,  1.33517,  1.33512,  1.33523,  1.33519,  1.33513,  1.33501,  1.33462,  1.33417,  1.33421,  1.33435,  1.33397,  1.33359,  1.33351,  1.33344,  1.33333,  1.33309,  1.33289,  1.33293,  1.33272,  1.33221,  1.33166,  1.33102,  1.33059,  1.33062,  1.33061,  1.33037,  1.33032,  1.33015,  1.32971,  1.32953,  1.32973,  1.32979,  1.32964,  1.32943,  1.32892,  1.32815,  1.32765,  1.32762,  1.32731,  1.32700,  1.32675,  1.32651,  1.32585,  1.32541,  1.32556,  1.32594,  1.32560,  1.32465,  1.32424,  1.32440,  1.32425,  1.32367,  1.32321,  1.32307,  1.32306,  1.32287,  1.32223,  1.32114,  1.32050,  1.32056,  1.32030,  1.31990,  1.31988,  1.31951,  1.31895,  1.31899,  1.31918,  1.31894,  1.31825,  1.31750,  1.31688,  1.31648,  1.31638,  1.31623,  1.31571,  1.31523,  1.31504,  1.31459,  1.31384,  1.31353,  1.31370,  1.31346,  1.31256,  1.31193,  1.31190,  1.31161,  1.31090,  1.31036,  1.31018,  1.31008,  1.30973,  1.30927,  1.30872,  1.30791,  1.30739,  1.30717,  1.30635,  1.30542,  1.30501,  1.30434,  1.30345,  1.30291,  1.30241,  1.30158,  1.30058,  1.29966,  1.29904,  1.29846,  1.29760,  1.29689,  1.29631,  1.29542,  1.29427,  1.29326,  1.29240,  1.29150,  1.29048,  1.28973,  1.28929,  1.28872,  1.28791,  1.28709,  1.28632,  1.28563,  1.28491,  1.28392,  1.28272,  1.28186,  1.28133,  1.28073,  1.27981,  1.27883,  1.27810,  1.27737,  1.27642,  1.27572,  1.27522,  1.27442,  1.27350,  1.27270,  1.27195,  1.27138,  1.27071,  1.26970,  1.26885,  1.26821,  1.26758,  1.26724,  1.26686,  1.26603,  1.26507,  1.26434,  1.26400,  1.26400,  1.26368,  1.26252,  1.26145,  1.26120,  1.26104,  1.26065,  1.26046,  1.26058,  1.26052,  1.25971,  1.25851,  1.25787,  1.25776,  1.25761,  1.25736,  1.25750,  1.25799,  1.25794,  1.25748,  1.25722,  1.25700,  1.25668,  1.25644,  1.25604,  1.25531,  1.25434,  1.25356,  1.25391,  1.25506,  1.25547,  1.25515,  1.25524,  1.25542,  1.25527,  1.25498,  1.25446,  1.25418,  1.25451,  1.25464,  1.25465,  1.25472,  1.25472,  1.25524,  1.25569,  1.25523,  1.25469,  1.25490,  1.25582,  1.25670,  1.25659,  1.25591,  1.25561,  1.25599,  1.25646,  1.25663,  1.25704,  1.25757,  1.25763,  1.25765,  1.25785,  1.25759,  1.25714,  1.25747,  1.25852,  1.25896,  1.25875,  1.25882,  1.25952,  1.26070,  1.26119,  1.26107,  1.26178,  1.26260,  1.26235,  1.26216,  1.26265,  1.26314,  1.26359,  1.26444,  1.26540,  1.26563,  1.26520,  1.26532,  1.26584,  1.26638,  1.26752,  1.26816,  1.26782,  1.26819,  1.26910,  1.26955,  1.26969,  1.26967,  1.27030,  1.27165,  1.27242,  1.27285,  1.27359,  1.27387,  1.27379,  1.27398,  1.27396,  1.27360,  1.27388,  1.27526,  1.27640,  1.27628,  1.27634,  1.27767,  1.27913,  1.27966,  1.27966,  1.27987,  1.28044,  1.28122,  1.28208,  1.28260,  1.28287,  1.28284,  1.28209,  1.28165,  1.28238,  1.28323,  1.28344,  1.28389,  1.28476,  1.28571,  1.28670,  1.28719,  1.28733,  1.28762,  1.28792,  1.28870,  1.28952,  1.28912,  1.28858,  1.28959,  1.29101,  1.29087,  1.28988,  1.28935,  1.28968,  1.29107,  1.29231,  1.29230,  1.29185,  1.29195,  1.29267,  1.29318,  1.29322,  1.29304,  1.29322,  1.29459,  1.29564,  1.29479,  1.29431,  1.29533,  1.29558,  1.29513,  1.29569,  1.29660,  1.29679,  1.29699,  1.29708,  1.29672,  1.29665,  1.29727,  1.29794,  1.29848,  1.29904,  1.29890,  1.29813,  1.29762,  1.29737,  1.29751,  1.29812,  1.29858,  1.29881,  1.29855,  1.29845,  1.29940,  1.30024,  1.30061,  1.30141,  1.30191,  1.30138,  1.30087,  1.30095,  1.30146,  1.30254,  1.30331,  1.30332,  1.30344,  1.30355,  1.30351,  1.30371,  1.30428,  1.30509,  1.30540,  1.30537,  1.30614,  1.30727,  1.30755,  1.30648,  1.30496,  1.30465,  1.30571,  1.30701,  1.30735,  1.30667,  1.30610,  1.30637,  1.30708,  1.30755,  1.30777,  1.30800,  1.30835,  1.30860,  1.30874,  1.30920,  1.30984,  1.31037,  1.31083,  1.31109,  1.31135,  1.31115,  1.31026,  1.31011,  1.31092,  1.31139,  1.31120,  1.31076,  1.31115,  1.31260,  1.31336,  1.31247,  1.31171,  1.31222,  1.31325,  1.31404,  1.31356,  1.31238,  1.31251,  1.31366,  1.31478,  1.31625,  1.31721,  1.31666,  1.31578,  1.31552,  1.31581,  1.31627,  1.31625,  1.31603,  1.31674,  1.31776,  1.31783,  1.31766,  1.31781,  1.31778,  1.31791,  1.31866,  1.31944,  1.31986,  1.32000,  1.32020,  1.32019,  1.31968,  1.31964,  1.32006,  1.32017,  1.32083,  1.32213,  1.32246,  1.32219,  1.32278,  1.32410,  1.32496,  1.32458,  1.32404,  1.32443,  1.32507,  1.32483,  1.32403,  1.32425,  1.32529,  1.32574,  1.32597,  1.32643,  1.32675,  1.32735,  1.32818,  1.32860,  1.32887,  1.32935,  1.33000,  1.33092,  1.33183,  1.33224,  1.33262,  1.33314,  1.33333,  1.33362,  1.33428,  1.33475,  1.33504,  1.33544,  1.33608,  1.33720,  1.33779,  1.33759,  1.33813,  1.33939,  1.34011,  1.34039,  1.34059,  1.34055,  1.34033,  1.33995,  1.34020,  1.34145,  1.34241,  1.34207,  1.34134,  1.34126,  1.34191,  1.34265,  1.34323,  1.34405,  1.34476,  1.34479,  1.34454,  1.34442,  1.34451,  1.34465,  1.34428,  1.34354,  1.34309,  1.34345,  1.34429,  1.34459,  1.34466,  1.34605,  1.34776,  1.34785,  1.34780,  1.34908,  1.35035,  1.35058,  1.35097,  1.35222,  1.35308,  1.35318,  1.35380,  1.35505,  1.35570,  1.35578,  1.35667,  1.35810,  1.35866,  1.35834,  1.35794,  1.35803,  1.35850,  1.35864,  1.35899,  1.36020,  1.36102,  1.36091,  1.36102,  1.36144,  1.36175,  1.36184,  1.36172,  1.36202,  1.36295,  1.36392,  1.36452,  1.36490,  1.36553,  1.36647,  1.36731,  1.36752,  1.36782,  1.36895,  1.36980,  1.37018,  1.37107,  1.37186,  1.37262,  1.37369,  1.37416,  1.37459,  1.37532,  1.37531,  1.37497,  1.37564,  1.37692,  1.37749,  1.37768,  1.37863,  1.37949,  1.37954,  1.37970,  1.37979,  1.37997,  1.38088,  1.38152,  1.38154,  1.38153,  1.38138,  1.38161,  1.38265,  1.38367,  1.38427,  1.38459,  1.38514,  1.38604,  1.38652,  1.38648,  1.38646,  1.38648,  1.38682,  1.38751,  1.38796,  1.38843,  1.38905,  1.38927,  1.38926,  1.38967,  1.39019,  1.39013,  1.38987,  1.39022,  1.39110,  1.39145,  1.39107,  1.39083,  1.39113,  1.39179,  1.39246,  1.39278,  1.39306,  1.39365,  1.39417,  1.39418,  1.39384,  1.39393,  1.39440,  1.39436,  1.39394,  1.39420,  1.39477,  1.39463,  1.39421,  1.39404,  1.39396,  1.39414,  1.39447,  1.39440,  1.39412,  1.39459,  1.39529,  1.39518,  1.39497,  1.39520,  1.39553,  1.39568,  1.39558,  1.39581,  1.39632,  1.39647,  1.39642,  1.39615,  1.39544,  1.39494,  1.39526,  1.39592,  1.39647,  1.39663,  1.39632,  1.39624,  1.39649,  1.39619,  1.39537,  1.39514,  1.39577,  1.39669,  1.39725,  1.39710,  1.39675,  1.39695,  1.39728,  1.39716,  1.39687,  1.39654,  1.39641,  1.39656,  1.39676,  1.39665,  1.39643,  1.39649,  1.39692,  1.39752,  1.39798,  1.39779,  1.39704,  1.39692,  1.39777,  1.39827,  1.39805,  1.39794,  1.39790,  1.39797,  1.39832,  1.39846,  1.39829,  1.39813,  1.39782,  1.39767,  1.39821,  1.39873,  1.39883,  1.39905,  1.39944,  1.39970,  1.39960,  1.39920,  1.39922,  1.39966,  1.40005,  1.40022,  1.40028,  1.40037,  1.40024,  1.39994,  1.40011,  1.40071,  1.40079,  1.40032,  1.40005,  1.40005,  1.40022,  1.40060,  1.40116,  1.40159,  1.40167,  1.40174,  1.40187,  1.40169,  1.40169,  1.40231,  1.40275,  1.40242,  1.40192,  1.40184,  1.40201,  1.40231,  1.40275,  1.40282,  1.40256,  1.40231,  1.40207,  1.40218,  1.40268,  1.40286,  1.40263,  1.40256,  1.40268,  1.40287,  1.40310,  1.40351,  1.40418,  1.40481,  1.40524,  1.40558,  1.40560,  1.40517,  1.40495,  1.40535,  1.40557,  1.40495,  1.40420,  1.40383,  1.40385,  1.40453,  1.40536,  1.40548,  1.40505,  1.40480,  1.40492,  1.40530,  1.40536,  1.40496,  1.40475,  1.40469,  1.40461,  1.40489,  1.40526,  1.40547,  1.40548,  1.40475,  1.40399,  1.40421,  1.40475,  1.40509,  1.40523,  1.40474,  1.40400,  1.40391,  1.40404,  1.40365,  1.40329,  1.40352,  1.40347,  1.40259,  1.40199,  1.40223,  1.40234,  1.40186,  1.40135,  1.40112,  1.40097,  1.40056,  1.39991,  1.39945,  1.39955,  1.39991,  1.39997,  1.39988,  1.39983,  1.39978,  1.39980,  1.39979,  1.39971,  1.39971,  1.39979,  1.39941,  1.39822,  1.39709,  1.39685,  1.39696,  1.39692,  1.39677,  1.39713,  1.39762,  1.39698,  1.39602,  1.39600,  1.39615,  1.39608,  1.39626,  1.39655,  1.39632,  1.39548,  1.39472,  1.39434,  1.39392,  1.39369,  1.39381,  1.39373,  1.39353,  1.39342,  1.39327,  1.39321,  1.39296,  1.39230,  1.39183,  1.39186,  1.39207,  1.39236,  1.39260,  1.39232,  1.39147,  1.39113,  1.39181,  1.39232,  1.39196,  1.39162,  1.39204,  1.39250,  1.39237,  1.39226,  1.39244,  1.39208,  1.39148,  1.39191,  1.39286,  1.39284,  1.39255,  1.39296,  1.39291,  1.39234,  1.39219,  1.39221,  1.39249,  1.39309,  1.39340,  1.39345,  1.39343,  1.39340,  1.39362,  1.39385,  1.39368,  1.39350,  1.39395,  1.39447,  1.39452,  1.39437,  1.39422,  1.39421,  1.39466,  1.39528,  1.39566,  1.39591,  1.39588,  1.39564,  1.39572,  1.39614,  1.39633,  1.39632,  1.39642,  1.39662,  1.39662,  1.39660,  1.39687,  1.39710,  1.39718,  1.39728,  1.39734,  1.39710,  1.39674,  1.39678,  1.39713,  1.39695,  1.39641,  1.39632,  1.39647,  1.39635,  1.39633,  1.39677,  1.39701,  1.39653,  1.39593,  1.39558,  1.39509,  1.39471,  1.39503,  1.39536,  1.39486,  1.39422,  1.39397,  1.39374,  1.39366,  1.39385,  1.39400,  1.39366,  1.39289,  1.39240,  1.39229,  1.39218,  1.39211,  1.39206,  1.39177,  1.39156,  1.39172,  1.39167,  1.39091,  1.38977,  1.38914,  1.38920,  1.38925,  1.38878,  1.38785,  1.38725,  1.38743,  1.38736,  1.38655,  1.38605,  1.38620,  1.38587,  1.38464,  1.38373,  1.38362,  1.38335,  1.38281,  1.38236,  1.38171,  1.38099,  1.38034,  1.37977,  1.37949,  1.37917,  1.37857,  1.37805,  1.37785,  1.37760,  1.37705,  1.37654,  1.37576,  1.37434,  1.37325,  1.37297,  1.37276,  1.37220,  1.37171,  1.37149,  1.37108,  1.37055,  1.37007,  1.36873,  1.36682,  1.36591,  1.36603,  1.36611,  1.36583,  1.36519,  1.36451,  1.36404,  1.36317,  1.36174,  1.36060,  1.36000,  1.35955,  1.35924,  1.35895,  1.35841,  1.35788,  1.35721,  1.35597,  1.35505,  1.35493,  1.35462,  1.35354,  1.35236,  1.35163,  1.35097,  1.34983,  1.34878,  1.34829,  1.34796,  1.34773,  1.34732,  1.34625,  1.34496,  1.34420,  1.34390,  1.34403,  1.34438,  1.34410,  1.34291,  1.34152,  1.34059,  1.33943,  1.33815,  1.33839,  1.33900,  1.33762,  1.33563,  1.33491,  1.33460,  1.33411,  1.33365,  1.33301,  1.33211,  1.33141,  1.33116,  1.33116,  1.33081,  1.32972,  1.32854,  1.32778,  1.32722,  1.32694,  1.32707,  1.32646,  1.32503,  1.32470,  1.32540,  1.32486,  1.32310,  1.32204,  1.32199,  1.32195,  1.32170,  1.32140,  1.32084,  1.32014,  1.31942,  1.31889,  1.31881,  1.31871,  1.31860,  1.31852,  1.31788,  1.31751,  1.31786,  1.31785,  1.31746,  1.31751,  1.31782,  1.31765,  1.31699,  1.31648,  1.31653,  1.31667,  1.31661,  1.31679,  1.31708,  1.31714,  1.31724,  1.31739,  1.31763,  1.31848,  1.31950,  1.31968,  1.31917,  1.31910,  1.31991,  1.32058,  1.32067,  1.32085,  1.32110,  1.32145,  1.32223,  1.32300,  1.32384,  1.32486,  1.32558,  1.32649,  1.32796,  1.32911,  1.32981,  1.33102,  1.33246,  1.33322,  1.33437,  1.33635,  1.33802,  1.33962,  1.34131,  1.34262,  1.34395,  1.34510,  1.34620,  1.34814,  1.35005,  1.35102,  1.35228,  1.35416,  1.35579,  1.35766,  1.36023,  1.36241,  1.36339,  1.36431,  1.36641,  1.36878,  1.37102,  1.37393,  1.37714,  1.37996,  1.38250,  1.38480,  1.38754,  1.39089,  1.39375,  1.39636,  1.39924,  1.40207,  1.40500,  1.40803,  1.41068,  1.41338,  1.41652,  1.41941,  1.42209,  1.42533,  1.42851,  1.43058,  1.43191,  1.43382,  1.43730,  1.44091,  1.44286,  1.44440,  1.44648,  1.44825,  1.44996,  1.45204,  1.45375,  1.45464,  1.45537,  1.45653,  1.45796,  1.45927,  1.46051,  1.46168,  1.46292,  1.46434,  1.46542,  1.46563,  1.46548,  1.46624,  1.46748,  1.46760,  1.46695,  1.46683,  1.46663,  1.46632,  1.46680,  1.46693,  1.46582,  1.46508,  1.46526,  1.46472,  1.46307,  1.46206,  1.46177,  1.46054,  1.45884,  1.45794,  1.45727,  1.45577,  1.45358,  1.45185,  1.45068,  1.44933,  1.44786,  1.44585,  1.44329,  1.44123,  1.43954,  1.43782,  1.43652,  1.43519,  1.43285,  1.42984,  1.42762,  1.42633,  1.42414,  1.42130,  1.41947,  1.41768,  1.41532,  1.41350,  1.41145,  1.40916,  1.40742,  1.40545,  1.40354,  1.40221,  1.40016,  1.39726,  1.39518,  1.39395,  1.39260,  1.39140,  1.39047,  1.38881,  1.38623,  1.38364,  1.38144,  1.37958,  1.37803,  1.37629,  1.37410,  1.37232,  1.37145,  1.37017,  1.36748,  1.36476,  1.36358,  1.36274,  1.36102,  1.35959,  1.35850,  1.35651,  1.35432,  1.35297,  1.35234,  1.35159,  1.34973,  1.34756,  1.34559,  1.34338,  1.34172,  1.34046,  1.33869,  1.33701,  1.33581,  1.33401,  1.33140,  1.32953,  1.32853,  1.32674,  1.32486,  1.32377,  1.32200,  1.31955,  1.31744,  1.31600,  1.31477,  1.31266,  1.31104,  1.31073,  1.30932,  1.30708,  1.30599,  1.30455,  1.30251,  1.30121,  1.29976,  1.29816,  1.29722,  1.29634,  1.29465,  1.29196,  1.28959,  1.28891,  1.28768,  1.28521,  1.28364,  1.28273,  1.28158,  1.27918,  1.27548,  1.27277,  1.27113,  1.26885,  1.26633,  1.26397,  1.26134,  1.25833,  1.25576,  1.25449,  1.25289,  1.24963,  1.24628,  1.24324,  1.23901,  1.23477,  1.23259,  1.23143,  1.22896,  1.22539,  1.22203,  1.21917,  1.21692,  1.21525,  1.21369,  1.21194,  1.21017,  1.20862,  1.20721,  1.20598,  1.20560,  1.20462,  1.20120,  1.19726,  1.19541,  1.19462,  1.19317,  1.19123,  1.18942,  1.18785,  1.18675,  1.18650,  1.18605,  1.18464,  1.18372,  1.18378,  1.18375,  1.18325,  1.18270,  1.18281,  1.18298,  1.18216,  1.18155,  1.18210,  1.18292,  1.18322,  1.18318,  1.18274,  1.18163,  1.18083,  1.18035,  1.17839,  1.17569,  1.17431,  1.17283,  1.17004,  1.16777,  1.16588,  1.16220,  1.15736,  1.15336,  1.14986,  1.14571,  1.14086,  1.13570,  1.13057,  1.12598,  1.12217,  1.11915,  1.11603,  1.11206,  1.10828,  1.10519,  1.10256,  1.09986,  1.09669,  1.09459,  1.09435,  1.09439,  1.09422,  1.09533,  1.09762,  1.09988,  1.10211,  1.10527,  1.11020,  1.11592,  1.12109,  1.12625,  1.13218,  1.13917,  1.14636,  1.15211,  1.15805,  1.16578,  1.17288,  1.17945,  1.18713,  1.19479,  1.20220,  1.21016,  1.21823,  1.22561,  1.23144,  1.23674,  1.24395,  1.25215,  1.25910,  1.26615,  1.27418,  1.28258,  1.29258,  1.30340,  1.31300,  1.32241,  1.33353,  1.34691,  1.36069,  1.37230,  1.38315,  1.39682,  1.41283,  1.42701,  1.43862,  1.45100,  1.46573,  1.48133,  1.49605,  1.50992,  1.52220,  1.53261,  1.54243,  1.54961,  1.55472,  1.56263,  1.57032,  1.57502,  1.58249,  1.58947,  1.58747,  1.58445,  1.59003,  1.59796,  1.60152,  1.59946,  1.59427,  1.59172,  1.59236,  1.59281,  1.59124,  1.58860,  1.58909,  1.59206,  1.59323,  1.59079,  1.58542,  1.58015,  1.57634,  1.57183,  1.56397,  1.55636,  1.55364,  1.54973,  1.54268,  1.54191,  1.54696,  1.55094,  1.55141,  1.55087,  1.55693,  1.57119,  1.58547,  1.59684,  1.60998,  1.62536,  1.64085,  1.65855,  1.67998,  1.70233,  1.72291,  1.74315,  1.76480,  1.78511,  1.80551,  1.82645,  1.84360,  1.85990,  1.87802,  1.89273,  1.90489,  1.91839,  1.92885,  1.93532,  1.94195,  1.94868,  1.95358,  1.95603,  1.95750,  1.96001,  1.96127,  1.95934,  1.95613,  1.95267,  1.94850,  1.94304,  1.93748,  1.93326,  1.92874,  1.92318,  1.91755,  1.91329,  1.91335,  1.91533,  1.91406,  1.91135,  1.90779,  1.90308,  1.89880,  1.89203,  1.88571,  1.88464,  1.88162,  1.87264,  1.86527,  1.86117,  1.85616,  1.84963,  1.84178,  1.83411,  1.82877,  1.82301,  1.81484,  1.80672,  1.79995,  1.79300,  1.78356,  1.77323,  1.76529,  1.75990,  1.75391,  1.74477,  1.73760,  1.73696,  1.73924,  1.74097,  1.74364,  1.74831,  1.75507,  1.76446,  1.77565,  1.78887,  1.80695,  1.82836,  1.84739,  1.86314,  1.87831,  1.89497,  1.91339,  1.93017,  1.94396,  1.95668,  1.96806,  1.97737,  1.98556,  1.99147,  1.99484,  1.99575,  1.99420,  1.99238,  1.99142,  1.98987,  1.98738,  1.98421,  1.98016,  1.97541,  1.96988,  1.96375,  1.95704,  1.94994,  1.94269,  1.93568,  1.92906,  1.92286,  1.91679,  1.91090,  1.90549,  1.90057,  1.89581,  1.89110,  1.88637,  1.88159,  1.87674,  
1.757,    1.741,    1.726,    1.701,    1.681,    1.663,    1.643,    1.613,    1.596,    1.551,    
1.512,    1.512,    1.542,    1.621,    1.741,    1.869,    1.939,    1.946,    1.926,    1.892,    
1.842,    1.823,    1.804,    1.782,    1.781,    1.848,    1.881,    1.918,    1.939,    1.930  ;

 idx_rfr_H2SO4_300K_PaW75_rl =
 1.930, 1.939, 1.918, 1.881, 1.848, 1.781, 1.782, 1.804, 1.823, 1.842, 1.892, 1.926, 1.946, 1.939, 1.869, 1.741, 1.621, 1.542, 1.512, 1.512, 1.551, 1.596, 1.613, 1.643, 1.663, 1.681, 1.701, 1.726, 1.741, 1.757, 1.796, 1.844, 1.869, 1.916, 1.911, 1.904, 1.842, 1.739, 1.676, 1.663, 1.678, 1.717, 1.756, 1.788, 1.807, 1.822, 1.849, 1.882, 1.947, 1.944, 1.907, 1.807, 1.702, 1.624, 1.589, 1.590, 1.626, 1.655, 1.669, 1.666, 1.643, 1.545, 1.479, 1.421, 1.320, 1.241, 1.179, 1.161, 1.151, 1.145, 1.144, 1.136, 1.133, 1.142, 1.173, 1.192, 1.222, 1.249, 1.272, 1.297, 1.308, 1.323, 1.331, 1.340, 1.351, 1.361, 1.368, 1.384, 1.399, 1.413, 1.422, 1.428, 1.434, 1.433, 1.430, 1.427, 1.420, 1.410, 1.392, 1.371, 1.361, 1.356, 1.350, 1.341, 1.337, 1.336, 1.336, 1.339, 1.342, 1.347, 1.353, 1.366, 1.379, 1.384, 1.386, 1.384, 1.386, 1.395, 1.397, 1.405, 1.399, 1.400, 1.398, 1.396, 1.395, 1.395, 1.395, 1.396, 1.396, 1.397, 1.394, 1.388, 1.370, 1.357, 1.341, 1.325, 1.306, 1.296, 1.294, 1.292, 1.288, 1.284, 1.277, 1.273, 1.272, 1.277, 1.279, 1.293, 1.308, 1.320, 1.332, 1.344, 1.352, 1.358, 1.362, 1.367, 1.370, 1.374, 1.377, 
1.380, 1.382, 1.384, 1.386, 1.388, 1.389, 1.391, 1.392, 
1.393, 1.394, 1.396, 1.397, 1.398, 1.398, 1.399, 1.400, 1.402, 1.403, 
1.403, 1.404, 1.405, 1.406, 1.406, 1.407, 1.408, 1.409, 1.410, 1.410, 
1.411, 1.411, 1.412, 1.413, 1.413, 1.415, 1.416, 1.416, 1.417, 1.418, 
1.419, 1.420, 1.421, 1.421, 1.422, 1.422, 1.423, 1.423, 1.424, 1.424, 
1.425, 1.425, 1.425, 1.426, 1.426, 1.427, 1.427, 1.427, 1.427, 1.427, 
1.427, 1.427, 1.427, 1.427, 1.427, 1.428, 1.431, 1.432, 1.438, 1.452  ;

 idx_rfr_H2SO4_300K_PaW75_img =
 2.00E-01, 2.26E-01, 3.00E-01, 3.20E-01, 3.29E-01, 2.90E-01, 2.57E-01, 2.40E-01, 2.35E-01, 2.38E-01, 2.61E-01, 2.99E-01, 3.62E-01, 4.57E-01, 5.54E-01, 5.94E-01, 5.64E-01, 4.79E-01, 3.52E-01, 2.99E-01, 2.21E-01, 1.91E-01, 1.83E-01, 1.73E-01, 1.71E-01, 1.65E-01, 1.60E-01, 1.57E-01, 1.57E-01, 1.58E-01, 1.68E-01, 1.94E-01, 2.16E-01, 3.13E-01, 3.41E-01, 3.86E-01, 4.64E-01, 4.63E-01, 4.10E-01, 3.51E-01, 3.01E-01, 2.75E-01, 2.71E-01, 2.77E-01, 2.82E-01, 2.92E-01, 3.11E-01, 3.38E-01, 4.53E-01, 5.38E-01, 6.37E-01, 7.08E-01, 7.11E-01, 6.68E-01, 6.12E-01, 5.60E-01, 5.40E-01, 5.56E-01, 5.90E-01, 6.34E-01, 6.81E-01, 7.55E-01, 7.61E-01, 7.58E-01, 7.19E-01, 6.63E-01, 5.93E-01, 5.47E-01, 5.13E-01, 4.45E-01, 3.97E-01, 3.51E-01, 3.23E-01, 2.62E-01, 2.11E-01, 1.95E-01, 1.73E-01, 1.58E-01, 1.43E-01, 1.43E-01, 1.37E-01, 1.30E-01, 1.26E-01, 1.22E-01, 1.21E-01, 1.22E-01, 1.23E-01, 1.25E-01, 1.30E-01, 1.38E-01, 1.44E-01, 1.52E-01, 1.64E-01, 1.75E-01, 1.84E-01, 1.91E-01, 2.03E-01, 2.15E-01, 2.25E-01, 2.20E-01, 2.12E-01, 2.09E-01, 2.06E-01, 1.94E-01, 1.82E-01, 1.71E-01, 1.60E-01, 1.51E-01, 1.44E-01, 1.35E-01, 1.28E-01, 1.18E-01, 1.16E-01, 1.17E-01, 1.21E-01, 1.19E-01, 1.13E-01, 1.09E-01, 1.10E-01, 1.17E-01, 1.21E-01, 1.24E-01, 1.26E-01, 1.27E-01, 1.27E-01, 1.27E-01, 1.27E-01, 1.28E-01, 1.30E-01, 1.36E-01, 1.43E-01, 1.53E-01, 1.61E-01, 1.59E-01, 1.59E-01, 1.50E-01, 1.31E-01, 1.09E-01, 9.90E-02, 9.30E-02, 8.60E-02, 8.20E-02, 7.30E-02, 5.60E-02, 5.20E-02, 2.30E-02, 1.90E-02, 6.00E-03, 0.00E+00, 0.00E+00, 0.00E+00, 3.76E-03, 2.97E-03, 2.41E-03, 2.09E-03, 1.86E-03, 1.67E-03, 1.54E-03, 1.43E-03, 
1.35E-03, 1.30E-03, 1.26E-03, 1.24E-03, 1.11E-03, 7.96E-04, 5.95E-04, 5.37E-04, 
4.86E-04, 4.24E-04, 3.61E-04, 3.14E-04, 2.72E-04, 2.34E-04, 2.02E-04, 1.76E-04, 1.55E-04, 1.38E-04, 
1.25E-04, 1.17E-04, 1.10E-04, 1.02E-04, 8.78E-05, 6.16E-05, 3.89E-05, 2.59E-05, 1.98E-05, 1.59E-05, 
1.27E-05, 1.05E-05, 8.93E-06, 7.75E-06, 6.94E-06, 5.63E-06, 4.95E-06, 4.05E-06, 2.46E-06, 1.84E-06, 
1.60E-06, 1.50E-06, 1.48E-06, 1.52E-06, 1.53E-06, 1.41E-06, 1.03E-06, 6.05E-07, 3.62E-07, 2.84E-07, 
2.33E-07, 2.02E-07, 1.83E-07, 1.58E-07, 1.24E-07, 9.98E-08, 8.79E-08, 8.46E-08, 8.39E-08, 8.20E-08, 
7.84E-08, 6.83E-08, 4.80E-08, 3.58E-08, 2.79E-08, 2.07E-08, 0.00E+00, 0.00E+00, 0.00E+00, 0.00E+00  ;

 idx_rfr_H2SO4_215K_75_HSL88_rl =
1.526, 1.512, 1.496, 1.484, 1.464, 1.456, 1.454, 1.454, 1.452, 1.452, 1.448, 1.443, 
1.432, 1.425, 1.411, 1.405, 1.390, 1.362, 1.319, 1.288, 1.292, 1.366, 1.383, 1.420, 
1.435, 1.427, 1.411, 1.376, 1.485, 1.485, 1.421, 1.235, 1.148, 1.220, 1.457, 1.753, 
1.767, 1.704, 1.791, 2.128, 2.094, 1.805, 1.823, 2.024, 1.808, 1.790, 1.739, 1.663, 
1.656, 1.692, 2.003, 2.207, 2.041, 1.895, 1.809, 1.942, 1.993 ;

 idx_rfr_H2SO4_215K_75_HSL88_img =
1.07e-8, 1.07e-8, 1.07e-8, 1.07e-8, 1.07e-8, 1.07e-8, 1.07e-8, 1.07e-8, 1.56e-8, 2.12e-8, 1.90e-7, 1.60e-6, 
1.06e-5, 1.46e-4, 5.85e-4, 0.00134, 0.00192, 0.00399, 0.00604, 0.0875,  0.144,   0.178,   0.179,   0.165, 
0.151,   0.156,   0.137,   0.195,   0.195,   0.147,   0.0841,  0.166,   0.461,   0.709,   0.840,   0.817, 
0.604,   0.557,   0.736,   0.465,   0.306,   0.210,   0.433,   0.199,   0.110,   0.112,   0.134,   0.163, 
0.181,   0.463,   0.616,   0.166,   0.0940,  0.0558,  0.146,   0.187,   0.0274 ;
}

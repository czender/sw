// ncgen -b -o $DATA/aca/idx_rfr_SAJ93.nc $HOME/idx_rfr/idx_rfr_SAJ93.cdl
// ncks -C -H -s %9.5f -v bnd,idx_rfr_afghan_dust_img,idx_rfr_afghan_dust_rl $DATA/aca/idx_rfr_SAJ93.nc

netcdf idx_rfr_SAJ93 {
dimensions:
	bnd=180;
variables:

	:RCS_Header = "$Id$";
	:history = "";
	:source="
Thu Jun 11 10:53:22 MDT 1998
Received afghan_dust, which is based on SAJ93. 
Afghan dust is less optically active than Saharan dust of Vol73 but more than dust_like or mineral_dust aerosols of DKS91.
The original data were 177 measurements of the indices of refraction from 0.34 to 25.0 microns.
I prepended three lines of mineral_dust properties onto the afghan_dust to cover the range 0.2--0.34 microns.
The mineral_dust data come from DKS91, as stored in /home/zender/dst/idx_rfr_dks91.nc
From 0.34--25.0 microns the afghan_dust data are true Afghan dust.
These indices are also shown graphically in STB98.";

	float bnd(bnd);
	bnd:long_name = "Band center wavelength";
	bnd:units = "micron";
	bnd:C_format = "%.5g";

	float idx_rfr_afghan_dust_rl(bnd);
	idx_rfr_afghan_dust_rl:long_name = "Afghan dust real index of refraction";
	idx_rfr_afghan_dust_rl:units = "";
	idx_rfr_afghan_dust_rl:C_format = "%.4g";

	float idx_rfr_afghan_dust_img(bnd);
	idx_rfr_afghan_dust_img:long_name = "Afghan dust imaginary index of refraction";
	idx_rfr_afghan_dust_img:units = "";
	idx_rfr_afghan_dust_img:C_format = "%.3g";

data:	

bnd =   0.2, 0.25, 0.3,
0.34483, 0.35714, 0.37037, 0.38462, 0.40000, 0.41667, 0.43478, 0.45455, 0.47619, 0.50000, 0.52632, 0.55556, 0.58824, 0.62500, 0.66667, 0.71429, 0.76923, 0.83333, 0.90909, 2.50000, 2.56410, 2.63158, 2.65957, 2.68817, 2.70270, 2.71739, 2.74725, 2.76243, 2.77778, 2.78940, 2.79330, 2.82486, 2.85714, 2.89017, 2.90698, 2.92398, 2.94118, 2.95858, 2.97619, 2.99401, 3.01205, 3.03030, 3.06748, 3.12500, 3.16456, 3.22581, 3.26797, 3.33333, 3.36700, 3.38983, 3.42466, 3.44828, 3.47222, 3.49650, 3.52113, 3.54610, 3.57143, 3.70370, 3.84615, 3.96825, 4.00000, 4.03226, 4.16667, 4.34783, 4.54545, 4.76190, 4.95050, 4.97512, 5.00000, 5.07614, 5.15464, 5.19481, 5.22193, 5.26316, 5.29101, 5.37634, 5.43478, 5.49451, 5.52486, 5.55556, 5.61798, 5.71429, 5.84795, 5.95238, 6.06061, 6.09756, 6.13497, 6.21118, 6.25000, 6.36943, 6.45161, 6.53595, 6.62252, 6.66667, 6.77966, 6.94444, 6.99301, 7.04225, 7.09220, 7.14286, 7.16846, 7.19424, 7.24638, 7.29927, 7.35294, 7.40741, 7.46269, 7.69231, 7.87402, 8.00000, 8.33333, 8.47458, 8.62069, 8.69565, 8.92857, 9.09091, 9.25926, 9.38967, 9.52381, 9.61539, 9.75610, 9.90099,10.00000,10.10101,10.41667,10.52632,10.63830,10.86957,11.11111,11.23596,11.36364,11.49425,11.76471,11.90476,12.04819,12.19512,12.34568,12.50000,12.82051,12.98701,13.15790,13.33333,13.51351,13.69863,13.88889,13.92758,13.98601,14.08451,14.28571,14.49275,14.70588,15.38461,15.62500,16.12903,16.39344,16.66667,16.94915,17.39130,17.85714,18.18182,18.51852,18.86792,19.23077,19.60784,20.00000,20.40816,20.83333,21.27660,21.50538,21.73913,22.22222,22.72727,23.25581,23.52941,23.80952,24.39024,25.00000;

idx_rfr_afghan_dust_rl = 1.5300, 1.5300, 1.5300,
1.5589,1.5592,1.5592,1.5595,1.5595,1.5597,1.5596,1.5598,1.5598,1.5599,1.5598,1.56  ,1.5598,1.56  ,1.5599,1.56  ,1.5598,1.5599,1.5598,1.5518,1.5501,1.5476,1.5461,1.5442,1.543 ,1.542 ,1.5412,1.5428,1.5437,1.5429,1.5427,1.5439,1.5456,1.5486,1.5506,1.5535,1.5558,1.5573,1.558 ,1.5587,1.5584,1.5582,1.5573,1.5561,1.555 ,1.5537,1.5522,1.55  ,1.55  ,1.5502,1.5517,1.5518,1.551 ,1.551 ,1.5514,1.5503,1.5496,1.5458,1.5426,1.5431,1.5421,1.5419,1.5375,1.5338,1.5293,1.5244,1.5203,1.5203,1.5204,1.5177,1.5147,1.5152,1.5143,1.5134,1.5125,1.5112,1.5086,1.507 ,1.5079,1.5088,1.5051,1.5007,1.4996,1.4987,1.4909,1.4937,1.497 ,1.5012,1.4998,1.4939,1.4906,1.4867,1.4797,1.4773,1.4834,1.5057,1.5127,1.5171,1.5153,1.5142,1.5108,1.5122,1.5178,1.5157,1.5101,1.5101,1.507 ,1.5001,1.4934,1.4879,1.4715,1.4711,1.4649,1.4626,1.4626,1.4746,1.4798,1.4825,1.4915,1.5161,1.5611,1.6058,1.6284,1.6465,1.6494,1.65  ,1.6441,1.6443,1.6378,1.6368,1.645 ,1.6621,1.6461,1.6335,1.6109,1.5892,1.5751,1.5771,1.5917,1.6002,1.6015,1.6065,1.6004,1.5929,1.5768,1.5871,1.5886,1.5882,1.5735,1.5816,1.5804,1.5509,1.5361,1.535 ,1.5173,1.5083,1.4885,1.4815,1.4641,1.4731,1.4787,1.5152,1.5345,1.5484,1.5114,1.5219,1.5594,1.6501,1.6725,1.7097,1.691 ,1.7337,1.7625,1.8011,1.7861,1.7982,1.7573;

idx_rfr_afghan_dust_img = 0.0700, 0.0300, 0.0250,
0.0035,0.0034,0.0034,0.0032,0.0032,0.0031,0.0031,0.0031,0.0031,0.0031,0.0031,0.003 ,0.0031,0.0032,0.0032,0.0033,0.0034,0.0036,0.0039,0.0056,0.0051,0.0054,0.006 ,0.0065,0.0075,0.0088,0.0129,0.0153,0.0145,0.0146,0.0155,0.0182,0.0208,0.0228,0.0237,0.0238,0.0225,0.0204,0.0192,0.0173,0.0157,0.0146,0.0132,0.011 ,0.0105,0.0095,0.0091,0.0099,0.0115,0.0107,0.0134,0.0102,0.0103,0.011 ,0.0092,0.0086,0.0083,0.0083,0.0093,0.0118,0.0104,0.0098,0.0105,0.0121,0.0139,0.0168,0.0203,0.0214,0.0205,0.0218,0.0232,0.0255,0.0246,0.0264,0.0271,0.0275,0.029 ,0.0317,0.0344,0.0321,0.0324,0.0368,0.0447,0.047 ,0.0494,0.058 ,0.0601,0.0556,0.0551,0.0562,0.0604,0.064 ,0.0687,0.0775,0.093 ,0.1077,0.1027,0.0967,0.0922,0.0903,0.0894,0.0961,0.0891,0.0825,0.0855,0.0838,0.0844,0.0882,0.0916,0.0957,0.1144,0.1297,0.1337,0.1444,0.1751,0.1984,0.2062,0.2264,0.2571,0.2833,0.2874,0.2814,0.2655,0.2436,0.1879,0.1797,0.1719,0.1619,0.1525,0.148 ,0.1647,0.1375,0.1054,0.0941,0.0834,0.0933,0.1106,0.1298,0.141 ,0.1388,0.1366,0.1306,0.121 ,0.119 ,0.1244,0.1325,0.1253,0.1149,0.1319,0.1338,0.1238,0.1236,0.1275,0.158 ,0.1468,0.1633,0.176 ,0.2081,0.2452,0.2783,0.3162,0.3404,0.3469,0.3348,0.3415,0.4239,0.4727,0.4976,0.4879,0.4516,0.4486,0.4654,0.4628,0.4426,0.4295,0.3943,0.4268;
}


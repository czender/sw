// $Id$
// ncgen -b -o ${DATA}/aca/idx_rfr_limestone.nc ${HOME}/idx_rfr/idx_rfr_limestone.cdl
// scp ${DATA}/aca/idx_rfr_limestone.nc ${HOME}/idx_rfr/idx_rfr_limestone.cdl dust.ess.uci.edu:/var/www/html/idx_rfr

netcdf idx_rfr_limestone {

dimensions:
	bnd_limestone_krk_QOL78 = 797 ;
variables:

// global attributes:
	:RCS_Header = "$Id$" ;
	:history = "" ;
	:description = "Refractive indices from QOL78" ;
	:source="
Charlie Zender (UCI) <zender at uci dot edu> created 20060619.

This file contains continuous refractive indices for
limstone from the UV to the IR.
Data from ~0.2--32.8 um comes from QOL78 as communicated by Ted Roush.
See also notes for limestone properties from QOL78 Lorentz dispersion method in idx_rfr.cc
Source file for QOL78 Kramers-Kronig data is Ted Roush in roush/limestone.oc.
Roush supplied an original e-mail with a naked table, and a processed
version of the table which he had annotated.
I attached the header from the latter to the table in the former
and converted to CDL format on 20060619.

Limestone samples are from Bethany Falls.
Limestone is primarily randomly oriented microcrystals of calcite, with 
dolomite and organic fossil material as secondary constituents.
Hence limestone is also known as amorphous calcite.
Separate measurements were made to facilitate two analysis techniques, 
Kramers-Kronig (KK) and Lorentz disperion (LD).
The refractive indices resulting show reasonable agreement from 0.2--25 um.
QOL78 found LD real and imginary indices higher than KK in 25--32.8 um.
Probably due to assumptions in KK analysis.
LD measurements are preferred in this region.

Limestone results may be reported in NOAA 76022603:
Holland, W.E., M.R. Querry, and R.M. Coveney, Jr. (1975), Measurements of spectral reflectance and optical constants of selected rock samples for application to remote sensing of soil moisture, NOAA Report 76022603: 78 pp.
which may be another name for
Holland, W.E., M.R. Querry, and R.M. Coveney, Jr., Measurements of spectral reflectance and optical constants of selected rock samples for application to remote sensing of soil moisture, Completion Report, U.S. Dept. of Commerce grant 04-4-158-27, available from National Technical Information Service, Springfield, VA 22151
There is also
Jordan, Ray E., Jr., Querry, Marvin R., Holland, Wayne E., Osbourn, Gordon C., and Coveney, Raymond M., Jr. (1975), Reflectance and complex refractive index of polycrystalline limestone, J. Opt. Soc. Am. A, vol. 65, page 1170.

Reference QOL78:
Querry, M.R, G.C. Osbourn, K. Lies, R. Jordon, R. Coveney, Jr. (1978), Complex refractive index of limestone in the visible and infrared, Appl. Opt., 17(3), 353-356.

************************************************************************
Begin Letter from Ted Roush, 20060619
************************************************************************
Hi Charlie,
I am attaching two files that I believe contain the Querry limestone data.
lmstn.con is the original file I got several years ago.  I thought it was in
unusual column format, so I read it and wrote the other file I am including
here (limestone, col 1= wavelength micron, wavenumber cm-1, n, k).

I can't provide any information regarding how the numbers in the original
file were actually generated.  I ASSUME they were derived via the dispersion
parameters listed in Querry's original paper.  I do have a couple of
programs that would take the oscillator parameters and create n's and k's.
If you are interested in my attempting that I am afraid my schedule would
prevent me from doing so for about a month.

I hope these help!
Ted

Dr. Ted L. Roush
NASA Ames Research Center
MS 245-3
Moffett Field, CA  94035-1000
************************************************************************
End Letter from Ted Roush, 20060619
************************************************************************

************************************************************************
Begin Procedure to create netCDF from Roush file roush/limestone.oc
************************************************************************
tbl2cdf ~/limestone.txt ~/limestone.nc
ncdump ~/limestone.nc > ~/limestone.cdl

ncks -v bnd ~/limestone.nc | m
ncks -u -v bnd_limestone,idx_rfr_illite_rl,idx_rfr_illite_img -s '%f, ' ~/limestone.nc | m
************************************************************************
End Procedure to create netCDF from Roush file roush/limestone.oc
************************************************************************
	";

// Begin contents of file:

	float bnd_limestone_krk_QOL78(bnd_limestone_krk_QOL78) ;
		bnd_limestone_krk_QOL78:units = "microns" ;
		bnd_limestone_krk_QOL78:longname = "Band center wavelength, Limestone" ;
		bnd_limestone_krk_QOL78:C_format = "%.5g" ;

	float wvn_limestone_krk_QOL78(bnd_limestone_krk_QOL78) ;
		wvn_limestone_krk_QOL78:units = "cm-1" ;
		wvn_limestone_krk_QOL78:longname = "Band center wavenumber, Limestone" ;
		wvn_limestone_krk_QOL78:C_format = "%.5g" ;

	float idx_rfr_limestone_krk_QOL78_rl(bnd_limestone_krk_QOL78) ;
		idx_rfr_limestone_krk_QOL78_rl:units = "" ;
		idx_rfr_limestone_krk_QOL78_rl:longname = "Limestone refractive index, real part " ;
		idx_rfr_limestone_krk_QOL78_rl:C_format = "%.4g" ;

	float idx_rfr_limestone_krk_QOL78_img(bnd_limestone_krk_QOL78) ;
		idx_rfr_limestone_krk_QOL78_img:units = "" ;
		idx_rfr_limestone_krk_QOL78_img:longname = "Limestone refractive index, imag part " ;
		idx_rfr_limestone_krk_QOL78_img:C_format = "%.3g" ;

// End contents limestone.txt file:

data:

 bnd_limestone_krk_QOL78 = 0.2, 0.21, 0.22, 0.23, 0.24, 0.25, 0.26, 0.27, 0.28, 0.29, 
    0.3, 0.31, 0.32, 0.33, 0.34, 0.35, 0.36, 0.37, 0.38, 0.39, 0.4, 0.41, 
    0.42, 0.43, 0.44, 0.45, 0.46, 0.47, 0.48, 0.49, 0.5, 0.51, 0.52, 0.53, 
    0.54, 0.55, 0.56, 0.57, 0.58, 0.59, 0.6, 0.61, 0.62, 0.63, 0.64, 0.65, 
    0.66, 0.67, 0.68, 0.69, 0.7, 0.71, 0.72, 0.73, 0.74, 0.75, 0.76, 0.77, 
    0.78, 0.79, 0.8, 0.81, 0.82, 0.83, 0.84, 0.85, 0.86, 0.87, 0.88, 0.89, 
    0.9, 0.91, 0.92, 0.93, 0.94, 0.95, 0.96, 0.97, 0.98, 0.99, 1, 1.01, 1.02, 
    1.03, 1.04, 1.05, 1.06, 1.07, 1.08, 1.09, 1.1, 1.11, 1.12, 1.13, 1.14, 
    1.15, 1.16, 1.17, 1.18, 1.19, 1.2, 1.21, 1.22, 1.23, 1.24, 1.25, 1.26, 
    1.27, 1.28, 1.29, 1.3, 1.31, 1.32, 1.33, 1.34, 1.35, 1.36, 1.37, 1.38, 
    1.39, 1.4, 1.41, 1.42, 1.43, 1.44, 1.45, 1.46, 1.47, 1.48, 1.49, 1.5, 
    1.51, 1.52, 1.53, 1.54, 1.55, 1.56, 1.57, 1.58, 1.59, 1.6, 1.61, 1.62, 
    1.63, 1.64, 1.65, 1.66, 1.67, 1.68, 1.69, 1.7, 1.71, 1.72, 1.73, 1.74, 
    1.75, 1.76, 1.77, 1.78, 1.79, 1.8, 1.81, 1.82, 1.83, 1.84, 1.85, 1.86, 
    1.87, 1.88, 1.89, 1.9, 1.91, 1.92, 1.93, 1.94, 1.95, 1.96, 1.97, 1.98, 
    1.99, 2, 2.05, 2.1, 2.15, 2.2, 2.25, 2.3, 2.35, 2.4, 2.45, 2.5, 2.55, 
    2.6, 2.65, 2.7, 2.75, 2.8, 2.85, 2.9, 2.95, 3, 3.05, 3.1, 3.15, 3.2, 
    3.25, 3.3, 3.35, 3.4, 3.45, 3.5, 3.55, 3.6, 3.65, 3.7, 3.75, 3.8, 3.85, 
    3.9, 3.95, 4, 4.05, 4.1, 4.15, 4.2, 4.25, 4.3, 4.35, 4.4, 4.45, 4.5, 
    4.55, 4.6, 4.65, 4.7, 4.75, 4.8, 4.85, 4.9, 4.95, 5, 5.05, 5.1, 5.15, 
    5.2, 5.25, 5.3, 5.35, 5.4, 5.45, 5.5, 5.55, 5.6, 5.65, 5.7, 5.75, 5.8, 
    5.85, 5.9, 5.95, 6, 6.05, 6.1, 6.15, 6.2, 6.25, 6.3, 6.35, 6.4, 6.45, 
    6.5, 6.55, 6.6, 6.65, 6.7, 6.75, 6.8, 6.85, 6.9, 6.95, 7, 7.05, 7.1, 
    7.15, 7.2, 7.25, 7.3, 7.35, 7.4, 7.45, 7.5, 7.55, 7.6, 7.65, 7.7, 7.75, 
    7.8, 7.85, 7.9, 7.95, 8, 8.05, 8.1, 8.15, 8.2, 8.25, 8.3, 8.35, 8.4, 
    8.45, 8.5, 8.55, 8.6, 8.65, 8.7, 8.75, 8.8, 8.85, 8.9, 8.95, 9, 9.05, 
    9.1, 9.15, 9.2, 9.25, 9.3, 9.35, 9.4, 9.45, 9.5, 9.55, 9.6, 9.65, 9.7, 
    9.75, 9.8, 9.85, 9.9, 9.95, 10, 10.05, 10.1, 10.15, 10.2, 10.25, 10.3, 
    10.35, 10.4, 10.45, 10.5, 10.55, 10.6, 10.65, 10.7, 10.75, 10.8, 10.85, 
    10.9, 10.95, 11, 11.05, 11.1, 11.15, 11.2, 11.25, 11.3, 11.35, 11.4, 
    11.45, 11.5, 11.55, 11.6, 11.65, 11.7, 11.75, 11.8, 11.85, 11.9, 11.95, 
    12, 12.05, 12.1, 12.15, 12.2, 12.25, 12.3, 12.35, 12.4, 12.45, 12.5, 
    12.55, 12.6, 12.65, 12.7, 12.75, 12.8, 12.85, 12.9, 12.95, 13, 13.05, 
    13.1, 13.15, 13.2, 13.25, 13.3, 13.35, 13.4, 13.45, 13.5, 13.55, 13.6, 
    13.65, 13.7, 13.75, 13.8, 13.85, 13.9, 13.95, 14, 14.05, 14.1, 14.15, 
    14.2, 14.25, 14.3, 14.35, 14.4, 14.45, 14.5, 14.55, 14.6, 14.65, 14.7, 
    14.75, 14.8, 14.85, 14.9, 14.95, 15, 15.05, 15.1, 15.15, 15.2, 15.25, 
    15.3, 15.35, 15.4, 15.45, 15.5, 15.55, 15.6, 15.65, 15.7, 15.75, 15.8, 
    15.85, 15.9, 15.95, 16, 16.05, 16.1, 16.15, 16.2, 16.25, 16.3, 16.35, 
    16.4, 16.45, 16.5, 16.55, 16.6, 16.65, 16.7, 16.75, 16.8, 16.85, 16.9, 
    16.95, 17, 17.05, 17.1, 17.15, 17.2, 17.25, 17.3, 17.35, 17.4, 17.45, 
    17.5, 17.55, 17.6, 17.65, 17.7, 17.75, 17.8, 17.85, 17.9, 17.95, 18, 
    18.05, 18.1, 18.15, 18.2, 18.25, 18.3, 18.35, 18.4, 18.45, 18.5, 18.55, 
    18.6, 18.65, 18.7, 18.75, 18.8, 18.85, 18.9, 18.95, 19, 19.05, 19.1, 
    19.15, 19.2, 19.25, 19.3, 19.35, 19.4, 19.45, 19.5, 19.55, 19.6, 19.65, 
    19.7, 19.75, 19.8, 19.85, 19.9, 19.95, 20, 20.05, 20.1, 20.15, 20.2, 
    20.25, 20.3, 20.35, 20.4, 20.45, 20.5, 20.55, 20.6, 20.65, 20.7, 20.75, 
    20.8, 20.85, 20.9, 20.95, 21, 21.05, 21.1, 21.15, 21.2, 21.25, 21.3, 
    21.35, 21.4, 21.45, 21.5, 21.55, 21.6, 21.65, 21.7, 21.75, 21.8, 21.85, 
    21.9, 21.95, 22, 22.05, 22.1, 22.15, 22.2, 22.25, 22.3, 22.35, 22.4, 
    22.45, 22.5, 22.55, 22.6, 22.65, 22.7, 22.75, 22.8, 22.85, 22.9, 22.95, 
    23, 23.05, 23.1, 23.15, 23.2, 23.25, 23.3, 23.35, 23.4, 23.45, 23.5, 
    23.55, 23.6, 23.65, 23.7, 23.75, 23.8, 23.85, 23.9, 23.95, 24, 24.05, 
    24.1, 24.15, 24.2, 24.25, 24.3, 24.35, 24.4, 24.45, 24.5, 24.55, 24.6, 
    24.65, 24.7, 24.75, 24.8, 24.85, 24.9, 24.95, 25, 25.05, 25.1, 25.15, 
    25.2, 25.25, 25.3, 25.35, 25.4, 25.45, 25.5, 25.55, 25.6, 25.65, 25.7, 
    25.75, 25.8, 25.85, 25.9, 25.95, 26, 26.05, 26.1, 26.15, 26.2, 26.25, 
    26.3, 26.35, 26.4, 26.45, 26.5, 26.55, 26.6, 26.65, 26.7, 26.75, 26.8, 
    26.85, 26.9, 26.95, 27, 27.05, 27.1, 27.15, 27.2, 27.25, 27.3, 27.35, 
    27.4, 27.45, 27.5, 27.55, 27.6, 27.65, 27.7, 27.75, 27.8, 27.85, 27.9, 
    27.95, 28, 28.05, 28.1, 28.15, 28.2, 28.25, 28.3, 28.35, 28.4, 28.45, 
    28.5, 28.55, 28.6, 28.65, 28.7, 28.75, 28.8, 28.85, 28.9, 28.95, 29, 
    29.05, 29.1, 29.15, 29.2, 29.25, 29.3, 29.35, 29.4, 29.45, 29.5, 29.55, 
    29.6, 29.65, 29.7, 29.75, 29.8, 29.85, 29.9, 29.95, 30, 30.05, 30.1, 
    30.15, 30.2, 30.25, 30.3, 30.35, 30.4, 30.45, 30.5, 30.55, 30.6, 30.65, 
    30.7, 30.75, 30.8, 30.85, 30.9, 30.95, 31, 31.05, 31.1, 31.15, 31.2, 
    31.25, 31.3, 31.35, 31.4, 31.45, 31.5, 31.55, 31.6, 31.65, 31.7, 31.75, 
    31.8, 31.85, 31.9, 31.95, 32, 32.05, 32.1, 32.15, 32.2, 32.25, 32.3, 
    32.35, 32.4, 32.45, 32.5, 32.55, 32.6, 32.65, 32.7, 32.75, 32.8 ;

 wvn_limestone_krk_QOL78 = 50000, 47619.1, 45454.5, 43478.3, 41666.7, 40000, 38461.5, 
    37037, 35714.3, 34482.8, 33333.3, 32258.1, 31250, 30303, 29411.8, 
    28571.4, 27777.8, 27027, 26315.8, 25641, 25000, 24390.2, 23809.5, 
    23255.8, 22727.3, 22222.2, 21739.1, 21276.6, 20833.3, 20408.2, 20000, 
    19607.8, 19230.8, 18867.9, 18518.5, 18181.8, 17857.1, 17543.9, 17241.4, 
    16949.2, 16666.7, 16393.4, 16129, 15873, 15625, 15384.6, 15151.5, 
    14925.4, 14705.9, 14492.8, 14285.7, 14084.5, 13888.9, 13698.6, 13513.5, 
    13333.3, 13157.9, 12987, 12820.5, 12658.2, 12500, 12345.7, 12195.1, 
    12048.2, 11904.8, 11764.7, 11627.9, 11494.3, 11363.6, 11236, 11111.1, 
    10989, 10869.6, 10752.7, 10638.3, 10526.32, 10416.67, 10309.28, 10204.08, 
    10101.01, 10000, 9900.99, 9803.92, 9708.74, 9615.38, 9523.81, 9433.96, 
    9345.79, 9259.26, 9174.31, 9090.91, 9009.01, 8928.57, 8849.56, 8771.93, 
    8695.65, 8620.69, 8547.01, 8474.58, 8403.36, 8333.33, 8264.46, 8196.72, 
    8130.08, 8064.52, 8000, 7936.51, 7874.02, 7812.5, 7751.94, 7692.31, 
    7633.59, 7575.76, 7518.8, 7462.69, 7407.41, 7352.94, 7299.27, 7246.38, 
    7194.24, 7142.86, 7092.2, 7042.25, 6993.01, 6944.44, 6896.55, 6849.31, 
    6802.72, 6756.76, 6711.41, 6666.67, 6622.52, 6578.95, 6535.95, 6493.51, 
    6451.61, 6410.26, 6369.43, 6329.11, 6289.31, 6250, 6211.18, 6172.84, 
    6134.97, 6097.56, 6060.61, 6024.1, 5988.02, 5952.38, 5917.16, 5882.35, 
    5847.95, 5813.95, 5780.35, 5747.13, 5714.29, 5681.82, 5649.72, 5617.98, 
    5586.59, 5555.56, 5524.86, 5494.51, 5464.48, 5434.78, 5405.41, 5376.34, 
    5347.59, 5319.15, 5291.01, 5263.16, 5235.6, 5208.33, 5181.35, 5154.64, 
    5128.21, 5102.04, 5076.14, 5050.5, 5025.13, 5000, 4878.05, 4761.9, 
    4651.16, 4545.45, 4444.44, 4347.83, 4255.32, 4166.67, 4081.63, 4000, 
    3921.57, 3846.15, 3773.58, 3703.7, 3636.36, 3571.43, 3508.77, 3448.28, 
    3389.83, 3333.33, 3278.69, 3225.81, 3174.6, 3125, 3076.92, 3030.3, 
    2985.07, 2941.18, 2898.55, 2857.14, 2816.9, 2777.78, 2739.73, 2702.7, 
    2666.67, 2631.58, 2597.4, 2564.1, 2531.65, 2500, 2469.14, 2439.02, 
    2409.64, 2380.95, 2352.94, 2325.58, 2298.85, 2272.73, 2247.19, 2222.22, 
    2197.8, 2173.91, 2150.54, 2127.66, 2105.26, 2083.33, 2061.86, 2040.82, 
    2020.2, 2000, 1980.2, 1960.78, 1941.75, 1923.08, 1904.76, 1886.79, 
    1869.16, 1851.85, 1834.86, 1818.18, 1801.8, 1785.71, 1769.91, 1754.39, 
    1739.13, 1724.14, 1709.4, 1694.92, 1680.67, 1666.67, 1652.89, 1639.34, 
    1626.02, 1612.9, 1600, 1587.3, 1574.8, 1562.5, 1550.39, 1538.46, 1526.72, 
    1515.15, 1503.76, 1492.54, 1481.48, 1470.59, 1459.85, 1449.28, 1438.85, 
    1428.57, 1418.44, 1408.45, 1398.6, 1388.89, 1379.31, 1369.86, 1360.54, 
    1351.35, 1342.28, 1333.33, 1324.5, 1315.79, 1307.19, 1298.7, 1290.32, 
    1282.05, 1273.89, 1265.82, 1257.86, 1250, 1242.24, 1234.57, 1226.99, 
    1219.51, 1212.12, 1204.82, 1197.6, 1190.48, 1183.43, 1176.47, 1169.59, 
    1162.79, 1156.07, 1149.43, 1142.86, 1136.36, 1129.94, 1123.6, 1117.32, 
    1111.11, 1104.97, 1098.9, 1092.9, 1086.96, 1081.08, 1075.27, 1069.52, 
    1063.83, 1058.2, 1052.63, 1047.12, 1041.67, 1036.27, 1030.93, 1025.64, 
    1020.41, 1015.23, 1010.1, 1005.025, 1000, 995.025, 990.099, 985.222, 
    980.392, 975.61, 970.874, 966.184, 961.539, 956.938, 952.381, 947.867, 
    943.396, 938.967, 934.579, 930.233, 925.926, 921.659, 917.431, 913.242, 
    909.091, 904.977, 900.901, 896.861, 892.857, 888.889, 884.956, 881.057, 
    877.193, 873.362, 869.565, 865.801, 862.069, 858.369, 854.701, 851.064, 
    847.458, 843.882, 840.336, 836.82, 833.333, 829.875, 826.446, 823.045, 
    819.672, 816.327, 813.008, 809.717, 806.452, 803.213, 800, 796.813, 
    793.651, 790.514, 787.402, 784.314, 781.25, 778.21, 775.194, 772.201, 
    769.231, 766.284, 763.359, 760.456, 757.576, 754.717, 751.88, 749.064, 
    746.269, 743.494, 740.741, 738.007, 735.294, 732.601, 729.927, 727.273, 
    724.638, 722.022, 719.424, 716.846, 714.286, 711.744, 709.22, 706.714, 
    704.225, 701.754, 699.301, 696.864, 694.444, 692.042, 689.655, 687.285, 
    684.932, 682.594, 680.272, 677.966, 675.676, 673.401, 671.141, 668.896, 
    666.667, 664.452, 662.252, 660.066, 657.895, 655.738, 653.595, 651.466, 
    649.351, 647.249, 645.161, 643.087, 641.026, 638.978, 636.943, 634.921, 
    632.911, 630.915, 628.931, 626.959, 625, 623.053, 621.118, 619.195, 
    617.284, 615.385, 613.497, 611.621, 609.756, 607.903, 606.061, 604.23, 
    602.41, 600.601, 598.802, 597.015, 595.238, 593.472, 591.716, 589.97, 
    588.235, 586.51, 584.795, 583.09, 581.395, 579.71, 578.035, 576.369, 
    574.713, 573.066, 571.429, 569.801, 568.182, 566.572, 564.972, 563.38, 
    561.798, 560.224, 558.659, 557.103, 555.556, 554.017, 552.486, 550.964, 
    549.451, 547.945, 546.448, 544.959, 543.478, 542.005, 540.541, 539.084, 
    537.634, 536.193, 534.759, 533.333, 531.915, 530.504, 529.101, 527.704, 
    526.316, 524.934, 523.56, 522.193, 520.833, 519.481, 518.135, 516.796, 
    515.464, 514.139, 512.82, 511.509, 510.204, 508.906, 507.614, 506.329, 
    505.051, 503.778, 502.513, 501.253, 500, 498.753, 497.512, 496.278, 
    495.049, 493.827, 492.611, 491.4, 490.196, 488.998, 487.805, 486.618, 
    485.437, 484.262, 483.092, 481.928, 480.769, 479.616, 478.469, 477.327, 
    476.19, 475.059, 473.934, 472.813, 471.698, 470.588, 469.484, 468.384, 
    467.29, 466.2, 465.116, 464.037, 462.963, 461.894, 460.829, 459.77, 
    458.716, 457.666, 456.621, 455.581, 454.545, 453.515, 452.489, 451.467, 
    450.45, 449.438, 448.431, 447.427, 446.429, 445.434, 444.444, 443.459, 
    442.478, 441.501, 440.529, 439.56, 438.596, 437.637, 436.681, 435.73, 
    434.783, 433.84, 432.9, 431.965, 431.034, 430.108, 429.185, 428.266, 
    427.35, 426.439, 425.532, 424.628, 423.729, 422.833, 421.941, 421.053, 
    420.168, 419.287, 418.41, 417.537, 416.667, 415.8, 414.938, 414.079, 
    413.223, 412.371, 411.523, 410.678, 409.836, 408.998, 408.163, 407.332, 
    406.504, 405.68, 404.858, 404.04, 403.226, 402.414, 401.606, 400.802, 
    400, 399.202, 398.406, 397.614, 396.825, 396.04, 395.257, 394.477, 
    393.701, 392.927, 392.157, 391.389, 390.625, 389.864, 389.105, 388.35, 
    387.597, 386.847, 386.1, 385.356, 384.615, 383.877, 383.142, 382.409, 
    381.679, 380.952, 380.228, 379.507, 378.788, 378.072, 377.358, 376.648, 
    375.94, 375.235, 374.532, 373.832, 373.134, 372.439, 371.747, 371.057, 
    370.37, 369.686, 369.004, 368.324, 367.647, 366.972, 366.3, 365.631, 
    364.964, 364.299, 363.636, 362.976, 362.319, 361.664, 361.011, 360.36, 
    359.712, 359.066, 358.423, 357.782, 357.143, 356.506, 355.872, 355.24, 
    354.61, 353.982, 353.357, 352.734, 352.113, 351.494, 350.877, 350.263, 
    349.65, 349.04, 348.432, 347.826, 347.222, 346.62, 346.021, 345.423, 
    344.828, 344.234, 343.643, 343.053, 342.466, 341.88, 341.297, 340.715, 
    340.136, 339.559, 338.983, 338.409, 337.838, 337.268, 336.7, 336.134, 
    335.57, 335.008, 334.448, 333.89, 333.333, 332.779, 332.226, 331.675, 
    331.126, 330.579, 330.033, 329.489, 328.947, 328.407, 327.869, 327.332, 
    326.797, 326.264, 325.733, 325.203, 324.675, 324.149, 323.625, 323.102, 
    322.581, 322.061, 321.543, 321.027, 320.513, 320, 319.489, 318.979, 
    318.471, 317.965, 317.46, 316.957, 316.456, 315.956, 315.457, 314.961, 
    314.465, 313.972, 313.48, 312.989, 312.5, 312.012, 311.526, 311.042, 
    310.559, 310.078, 309.598, 309.119, 308.642, 308.166, 307.692, 307.22, 
    306.748, 306.279, 305.81, 305.344, 304.878 ;

 idx_rfr_limestone_krk_QOL78_rl = 
	// CSZ 20060620: 
	// Values at 0.20 um are anomalous due to Kramers-Kronig boundary condition
	// Replace values at 0.20 um with values at 0.21 um
//	1.277, 
    1.613, 
    1.613, 1.6, 1.592, 1.584, 1.583, 1.593, 1.588, 
    1.579, 1.579, 1.569, 1.564, 1.563, 1.559, 1.554, 1.553, 1.551, 1.55, 
    1.548, 1.549, 1.548, 1.549, 1.557, 1.566, 1.57, 1.571, 1.566, 1.568, 
    1.569, 1.569, 1.566, 1.561, 1.561, 1.562, 1.562, 1.562, 1.562, 1.561, 
    1.562, 1.561, 1.565, 1.569, 1.568, 1.567, 1.569, 1.568, 1.567, 1.563, 
    1.56, 1.56, 1.556, 1.551, 1.55, 1.549, 1.552, 1.549, 1.55, 1.551, 1.552, 
    1.551, 1.552, 1.552, 1.555, 1.55, 1.55, 1.552, 1.552, 1.554, 1.555, 
    1.555, 1.554, 1.551, 1.553, 1.555, 1.555, 1.557, 1.56, 1.559, 1.56, 1.56, 
    1.562, 1.564, 1.564, 1.564, 1.562, 1.564, 1.564, 1.564, 1.563, 1.564, 
    1.563, 1.563, 1.564, 1.568, 1.565, 1.563, 1.565, 1.564, 1.563, 1.564, 
    1.564, 1.565, 1.564, 1.565, 1.566, 1.566, 1.566, 1.566, 1.567, 1.567, 
    1.566, 1.566, 1.568, 1.568, 1.568, 1.567, 1.566, 1.567, 1.567, 1.567, 
    1.567, 1.567, 1.567, 1.567, 1.567, 1.567, 1.568, 1.568, 1.568, 1.568, 
    1.568, 1.568, 1.568, 1.569, 1.569, 1.569, 1.569, 1.568, 1.568, 1.569, 
    1.568, 1.569, 1.568, 1.569, 1.568, 1.569, 1.568, 1.569, 1.569, 1.569, 
    1.569, 1.569, 1.568, 1.569, 1.567, 1.569, 1.568, 1.569, 1.57, 1.569, 
    1.569, 1.568, 1.568, 1.567, 1.567, 1.566, 1.565, 1.565, 1.564, 1.563, 
    1.563, 1.563, 1.563, 1.563, 1.563, 1.564, 1.563, 1.563, 1.563, 1.565, 
    1.571, 1.582, 1.581, 1.579, 1.579, 1.576, 1.571, 1.568, 1.575, 1.572, 
    1.566, 1.573, 1.586, 1.575, 1.623, 1.638, 1.511, 1.476, 1.51, 1.527, 
    1.535, 1.546, 1.543, 1.535, 1.541, 1.542, 1.536, 1.532, 1.531, 1.53, 
    1.534, 1.532, 1.532, 1.531, 1.528, 1.523, 1.519, 1.516, 1.513, 1.508, 
    1.518, 1.511, 1.507, 1.503, 1.502, 1.492, 1.467, 1.491, 1.489, 1.483, 
    1.481, 1.48, 1.476, 1.471, 1.468, 1.466, 1.462, 1.457, 1.451, 1.446, 
    1.441, 1.436, 1.423, 1.412, 1.406, 1.4, 1.393, 1.387, 1.377, 1.365, 
    1.347, 1.327, 1.352, 1.332, 1.316, 1.302, 1.286, 1.267, 1.242, 1.217, 
    1.188, 1.167, 1.127, 1.087, 1.038, 0.987, 0.895, 0.816, 0.646, 0.421, 
    0.403, 0.476, 0.543, 0.633, 0.74, 0.871, 1.036, 1.251, 1.47, 1.731, 
    2.016, 2.481, 2.91, 2.977, 2.762, 2.581, 2.424, 2.312, 2.23, 2.175, 
    2.114, 2.079, 2.034, 2.002, 1.979, 1.946, 1.923, 1.902, 1.877, 1.862, 
    1.86, 1.858, 1.847, 1.832, 1.819, 1.811, 1.8, 1.794, 1.783, 1.781, 1.775, 
    1.768, 1.762, 1.758, 1.755, 1.747, 1.75, 1.743, 1.734, 1.736, 1.732, 
    1.731, 1.723, 1.72, 1.723, 1.717, 1.717, 1.716, 1.715, 1.708, 1.703, 
    1.703, 1.698, 1.694, 1.702, 1.696, 1.688, 1.684, 1.687, 1.684, 1.681, 
    1.678, 1.675, 1.672, 1.664, 1.661, 1.656, 1.651, 1.643, 1.637, 1.627, 
    1.622, 1.613, 1.604, 1.596, 1.586, 1.576, 1.562, 1.545, 1.522, 1.497, 
    1.46, 1.403, 1.328, 1.242, 1.191, 1.246, 1.46, 1.844, 2.237, 2.286, 
    2.123, 1.971, 1.895, 1.83, 1.795, 1.775, 1.761, 1.743, 1.729, 1.713, 
    1.707, 1.697, 1.691, 1.683, 1.68, 1.675, 1.67, 1.671, 1.661, 1.66, 1.656, 
    1.65, 1.645, 1.64, 1.636, 1.632, 1.63, 1.624, 1.621, 1.617, 1.61, 1.608, 
    1.608, 1.6, 1.596, 1.589, 1.587, 1.58, 1.577, 1.571, 1.564, 1.557, 1.547, 
    1.537, 1.524, 1.505, 1.475, 1.431, 1.417, 1.485, 1.608, 1.673, 1.651, 
    1.622, 1.605, 1.592, 1.582, 1.575, 1.569, 1.566, 1.561, 1.555, 1.554, 
    1.548, 1.543, 1.538, 1.535, 1.537, 1.529, 1.516, 1.516, 1.516, 1.514, 
    1.512, 1.509, 1.508, 1.504, 1.5, 1.497, 1.494, 1.494, 1.491, 1.489, 
    1.486, 1.484, 1.481, 1.479, 1.476, 1.475, 1.472, 1.47, 1.466, 1.464, 
    1.463, 1.458, 1.457, 1.455, 1.451, 1.452, 1.447, 1.446, 1.444, 1.442, 
    1.439, 1.436, 1.434, 1.433, 1.43, 1.424, 1.425, 1.424, 1.423, 1.422, 
    1.421, 1.418, 1.416, 1.414, 1.409, 1.409, 1.407, 1.403, 1.399, 1.399, 
    1.393, 1.391, 1.388, 1.386, 1.383, 1.38, 1.377, 1.372, 1.37, 1.368, 
    1.366, 1.364, 1.358, 1.355, 1.352, 1.35, 1.348, 1.343, 1.339, 1.338, 
    1.334, 1.334, 1.329, 1.324, 1.324, 1.322, 1.318, 1.312, 1.308, 1.308, 
    1.307, 1.3, 1.298, 1.296, 1.291, 1.288, 1.286, 1.28, 1.277, 1.278, 1.272, 
    1.271, 1.264, 1.258, 1.257, 1.253, 1.249, 1.242, 1.238, 1.236, 1.232, 
    1.229, 1.222, 1.218, 1.214, 1.211, 1.208, 1.202, 1.197, 1.195, 1.192, 
    1.189, 1.183, 1.179, 1.179, 1.174, 1.173, 1.17, 1.167, 1.17, 1.168, 
    1.164, 1.159, 1.157, 1.157, 1.154, 1.151, 1.145, 1.141, 1.141, 1.138, 
    1.136, 1.129, 1.125, 1.122, 1.117, 1.112, 1.104, 1.099, 1.096, 1.091, 
    1.085, 1.078, 1.072, 1.069, 1.064, 1.058, 1.049, 1.042, 1.038, 1.032, 
    1.026, 1.016, 1.009, 1.005, 0.998, 0.992, 0.982, 0.976, 0.972, 0.965, 
    0.959, 0.95, 0.943, 0.939, 0.932, 0.926, 0.917, 0.91, 0.905, 0.897, 
    0.891, 0.88, 0.866, 0.853, 0.847, 0.845, 0.838, 0.83, 0.823, 0.813, 
    0.803, 0.792, 0.781, 0.772, 0.761, 0.751, 0.739, 0.728, 0.716, 0.705, 
    0.695, 0.685, 0.678, 0.668, 0.658, 0.647, 0.62, 0.601, 0.594, 0.56, 
    0.554, 0.545, 0.532, 0.521, 0.512, 0.5, 0.49, 0.479, 0.466, 0.456, 0.443, 
    0.435, 0.427, 0.408, 0.387, 0.365, 0.353, 0.343, 0.337, 0.331, 0.323, 
    0.315, 0.31, 0.299, 0.3, 0.295, 0.293, 0.271, 0.255, 0.245, 0.246, 0.247, 
    0.247, 0.243, 0.239, 0.233, 0.226, 0.225, 0.216, 0.216, 0.213, 0.213, 
    0.211, 0.208, 0.205, 0.201, 0.2, 0.2, 0.194, 0.192, 0.189, 0.193, 0.19, 
    0.185, 0.193, 0.189, 0.184, 0.176, 0.175, 0.172, 0.158, 0.169, 0.158, 
    0.146, 0.165, 0.136, 0.174, 0.147, 0.145, 0.156, 0.157, 0.163, 0.165, 
    0.155, 0.162, 0.159, 0.164, 0.165, 0.159, 0.158, 0.158, 0.156, 0.158, 
    0.152, 0.159, 0.156, 0.161, 0.162, 0.16, 0.156, 0.159, 0.163, 0.158, 
    0.141, 0.159, 0.149, 0.158, 0.158, 0.154, 0.158, 0.152, 0.174, 0.166, 
    0.165, 0.166, 0.175, 0.155, 0.136, 0.184, 0.207, 0.191, 0.154, 0.163, 
    0.156, 0.156, 0.191, 0.19, 0.192, 0.189, 0.189, 0.194, 0.203, 0.205, 
    0.201, 0.207, 0.205, 0.219, 0.229, 0.222, 0.229, 0.219, 0.258, 0.252, 
    0.252, 0.245, 0.255, 0.27, 0.276, 0.265, 0.28, 0.281, 0.307, 0.326, 
    0.323, 0.331, 0.324, 0.354, 0.357, 0.355, 0.355, 0.377, 
	// CSZ 20060620: 
	// Values at 32.8 um are anomalous due to Kramers-Kronig boundary condition
	// Replace values at 32.8 um with values at 32.75 um
	// 0.159 ;
	0.377 ; 

 idx_rfr_limestone_krk_QOL78_img = 
	// CSZ 20060620: 
	// Values at 0.20 um are anomalous due to Kramers-Kronig boundary condition
	// Replace values at 0.20 um with values at 0.21 um
	//	0.472, 
    0.058, 
    0.058, 0.052, 0.052, 0.054, 0.061, 0.055, 
    0.042, 0.041, 0.038, 0.034, 0.037, 0.037, 0.036, 0.037, 0.04, 0.042, 
    0.044, 0.047, 0.05, 0.052, 0.058, 0.064, 0.061, 0.055, 0.048, 0.047, 
    0.048, 0.044, 0.041, 0.037, 0.038, 0.041, 0.041, 0.04, 0.041, 0.04, 
    0.041, 0.041, 0.043, 0.045, 0.041, 0.038, 0.038, 0.036, 0.032, 0.029, 
    0.027, 0.028, 0.027, 0.025, 0.028, 0.032, 0.034, 0.035, 0.035, 0.038, 
    0.04, 0.04, 0.04, 0.041, 0.042, 0.04, 0.039, 0.044, 0.045, 0.046, 0.047, 
    0.046, 0.045, 0.044, 0.046, 0.049, 0.05, 0.051, 0.052, 0.051, 0.05, 0.05, 
    0.051, 0.052, 0.05, 0.049, 0.048, 0.049, 0.049, 0.048, 0.048, 0.048, 
    0.048, 0.047, 0.049, 0.051, 0.048, 0.045, 0.048, 0.048, 0.047, 0.048, 
    0.049, 0.049, 0.048, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.048, 0.049, 0.05, 0.048, 0.047, 0.047, 0.048, 0.048, 0.048, 
    0.048, 0.049, 0.049, 0.049, 0.049, 0.049, 0.05, 0.05, 0.049, 0.049, 0.05, 
    0.05, 0.049, 0.05, 0.05, 0.05, 0.049, 0.049, 0.049, 0.05, 0.049, 0.049, 
    0.05, 0.05, 0.049, 0.049, 0.05, 0.049, 0.05, 0.05, 0.05, 0.049, 0.049, 
    0.049, 0.05, 0.05, 0.051, 0.05, 0.051, 0.05, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.05, 0.05, 0.05, 0.051, 0.053, 0.054, 0.055, 0.056, 
    0.057, 0.058, 0.059, 0.06, 0.063, 0.068, 0.07, 0.059, 0.053, 0.05, 0.048, 
    0.045, 0.044, 0.049, 0.051, 0.045, 0.05, 0.058, 0.049, 0.06, 0.049, 
    0.049, 0.049, 0.018, 0.064, 0.073, 0.066, 0.061, 0.05, 0.05, 0.054, 
    0.049, 0.045, 0.05, 0.054, 0.057, 0.057, 0.055, 0.056, 0.054, 0.051, 
    0.05, 0.052, 0.054, 0.055, 0.061, 0.061, 0.053, 0.055, 0.055, 0.054, 
    0.044, 0.062, 0.078, 0.064, 0.066, 0.068, 0.067, 0.065, 0.066, 0.068, 
    0.067, 0.066, 0.065, 0.064, 0.064, 0.064, 0.06, 0.057, 0.062, 0.066, 
    0.068, 0.07, 0.069, 0.067, 0.067, 0.067, 0.089, 0.095, 0.072, 0.077, 
    0.075, 0.075, 0.071, 0.071, 0.074, 0.078, 0.084, 0.077, 0.085, 0.087, 
    0.096, 0.092, 0.147, 0.118, 0.357, 0.645, 0.856, 1.028, 1.191, 1.347, 
    1.49, 1.648, 1.747, 1.843, 1.871, 1.931, 1.867, 1.476, 0.912, 0.559, 
    0.408, 0.315, 0.282, 0.263, 0.243, 0.228, 0.219, 0.205, 0.207, 0.198, 
    0.191, 0.193, 0.189, 0.193, 0.205, 0.211, 0.203, 0.194, 0.192, 0.192, 
    0.192, 0.192, 0.193, 0.195, 0.198, 0.195, 0.195, 0.197, 0.199, 0.198, 
    0.199, 0.2, 0.193, 0.199, 0.201, 0.199, 0.198, 0.196, 0.202, 0.201, 
    0.199, 0.2, 0.199, 0.196, 0.193, 0.195, 0.194, 0.192, 0.199, 0.198, 
    0.188, 0.188, 0.191, 0.193, 0.189, 0.187, 0.184, 0.182, 0.179, 0.178, 
    0.177, 0.174, 0.172, 0.17, 0.169, 0.169, 0.169, 0.169, 0.171, 0.171, 
    0.171, 0.17, 0.17, 0.169, 0.17, 0.174, 0.176, 0.19, 0.233, 0.33, 0.507, 
    0.748, 0.977, 1.061, 0.819, 0.407, 0.185, 0.132, 0.128, 0.124, 0.14, 
    0.145, 0.145, 0.144, 0.145, 0.148, 0.152, 0.152, 0.155, 0.157, 0.159, 
    0.158, 0.161, 0.159, 0.156, 0.159, 0.155, 0.153, 0.154, 0.154, 0.154, 
    0.154, 0.154, 0.153, 0.153, 0.15, 0.151, 0.154, 0.151, 0.148, 0.149, 
    0.149, 0.15, 0.148, 0.149, 0.147, 0.147, 0.145, 0.145, 0.145, 0.145, 
    0.146, 0.154, 0.19, 0.274, 0.364, 0.368, 0.279, 0.208, 0.188, 0.179, 
    0.174, 0.173, 0.173, 0.172, 0.172, 0.169, 0.17, 0.169, 0.166, 0.167, 
    0.167, 0.169, 0.167, 0.16, 0.164, 0.172, 0.173, 0.173, 0.173, 0.174, 
    0.173, 0.172, 0.173, 0.174, 0.176, 0.178, 0.176, 0.177, 0.177, 0.178, 
    0.178, 0.179, 0.179, 0.18, 0.179, 0.18, 0.18, 0.18, 0.18, 0.18, 0.184, 
    0.182, 0.183, 0.183, 0.182, 0.186, 0.185, 0.184, 0.183, 0.184, 0.187, 
    0.186, 0.183, 0.186, 0.189, 0.191, 0.19, 0.187, 0.186, 0.186, 0.188, 
    0.185, 0.183, 0.185, 0.182, 0.184, 0.184, 0.181, 0.179, 0.182, 0.183, 
    0.183, 0.18, 0.18, 0.179, 0.182, 0.183, 0.18, 0.181, 0.179, 0.181, 0.181, 
    0.179, 0.181, 0.179, 0.181, 0.182, 0.18, 0.181, 0.181, 0.182, 0.182, 
    0.181, 0.179, 0.178, 0.181, 0.182, 0.181, 0.179, 0.178, 0.184, 0.18, 
    0.178, 0.18, 0.179, 0.182, 0.183, 0.18, 0.177, 0.178, 0.177, 0.177, 
    0.176, 0.174, 0.174, 0.176, 0.177, 0.174, 0.175, 0.174, 0.177, 0.177, 
    0.175, 0.177, 0.178, 0.18, 0.181, 0.18, 0.181, 0.181, 0.185, 0.185, 
    0.185, 0.185, 0.189, 0.191, 0.191, 0.19, 0.186, 0.186, 0.187, 0.186, 
    0.183, 0.181, 0.179, 0.18, 0.178, 0.176, 0.173, 0.171, 0.169, 0.166, 
    0.162, 0.161, 0.158, 0.159, 0.157, 0.154, 0.152, 0.151, 0.151, 0.149, 
    0.147, 0.144, 0.144, 0.142, 0.14, 0.139, 0.138, 0.137, 0.136, 0.135, 
    0.135, 0.135, 0.134, 0.134, 0.134, 0.133, 0.133, 0.133, 0.131, 0.131, 
    0.131, 0.131, 0.131, 0.127, 0.127, 0.126, 0.125, 0.123, 0.117, 0.114, 
    0.121, 0.128, 0.129, 0.124, 0.123, 0.122, 0.12, 0.12, 0.117, 0.117, 
    0.119, 0.119, 0.119, 0.118, 0.119, 0.121, 0.124, 0.127, 0.128, 0.129, 
    0.128, 0.128, 0.119, 0.115, 0.13, 0.125, 0.134, 0.153, 0.159, 0.166, 
    0.174, 0.18, 0.185, 0.195, 0.2, 0.206, 0.212, 0.219, 0.232, 0.233, 0.23, 
    0.237, 0.252, 0.277, 0.295, 0.306, 0.318, 0.327, 0.348, 0.359, 0.368, 
    0.379, 0.387, 0.396, 0.402, 0.414, 0.435, 0.453, 0.476, 0.487, 0.489, 
    0.497, 0.504, 0.528, 0.54, 0.544, 0.557, 0.566, 0.589, 0.6, 0.601, 0.608, 
    0.617, 0.643, 0.651, 0.651, 0.66, 0.67, 0.695, 0.701, 0.704, 0.711, 0.71, 
    0.73, 0.742, 0.742, 0.742, 0.758, 0.786, 0.785, 0.802, 0.799, 0.82, 
    0.848, 0.841, 0.857, 0.866, 0.871, 0.899, 0.9, 0.897, 0.906, 0.91, 0.939, 
    0.942, 0.934, 0.942, 0.946, 0.977, 0.986, 0.982, 0.988, 0.993, 1.025, 
    1.03, 1.018, 1.026, 1.033, 1.06, 1.059, 1.063, 1.073, 1.075, 1.113, 
    1.116, 1.11, 1.114, 1.128, 1.159, 1.157, 1.149, 1.158, 1.153, 1.175, 
    1.221, 1.228, 1.2, 1.168, 1.214, 1.241, 1.23, 1.26, 1.263, 1.284, 1.292, 
    1.276, 1.284, 1.291, 1.327, 1.331, 1.319, 1.324, 1.33, 1.375, 1.374, 
    1.359, 1.358, 1.378, 1.416, 1.408, 1.389, 1.397, 1.407, 1.445, 1.443, 
    1.432, 1.44, 1.445, 1.492, 1.485, 1.46, 1.452, 1.459, 1.496, 1.491, 
    1.466, 1.474, 1.477, 
	// CSZ 20060620: 
	// Values at 32.8 um are anomalous due to Kramers-Kronig boundary condition
	// Replace values at 32.8 um with values at 32.75 um
	// 0.031 ;
	1.477 ;

}

// $Id$
// ncgen -b -o ${DATA}/aca/idx_rfr_Ill_Kao_Mnt.nc ${HOME}/idx_rfr/idx_rfr_Ill_Kao_Mnt.cdl
// scp ${DATA}/aca/idx_rfr_Ill_Kao_Mnt.nc ${HOME}/idx_rfr/idx_rfr_Ill_Kao_Mnt.cdl dust.ess.uci.edu:/var/www/html/idx_rfr

netcdf idx_rfr_Ill_Kao_Mnt {

dimensions:
//	bnd_illite = 44 ;
	bnd_illite = 3994 ;
	bnd_kaolinite = 3994 ;
	bnd_montmorillonite = 444 ;
variables:

// global attributes:
	:RCS_Header = "$Id$" ;
	:history = "" ;
	:description = "Merged refractive indices from EgH79 and Roush" ;
	:source="
Charlie Zender (UCI) <zender at uci dot edu> created 20060512.

This file contains best-guess continuous refractive indices for
Illite, Kaolinite, and Montmorillonite from the UV to the IR.
In all cases the data from ~0.2--2.5 um comes from EgH79,
and the NIR--IR data come from Roush.
The mid-infrared Illite data were measured by Marvin Querry and reported in 1987 
U.S. Army tech. note CRDEC-CR-88009 from Aberdeen, MD.
The mid-infrared Kaolinite and Montmorillonite data were measured by Roush
and reported in RPO91.

The source files are idx_rfr_EgH79.nc and idx_rfr_roush_*.nc.
Roush supplied two flavors of Kaolinite, named kaolinite_1 and kaolinite_2.
I chose kaolinite_2 for this merged file since kaolinite_2 has 
has wider range and higher resolution (1 cm-1) than kaolinite_1.

Roush supplied two flavors of Montmorillonite, named montmorillonite_1
(from Clay Spur, Wyoming), and montmorillonite_2 (from Amory, Mississippi), 
respectively. 
I rather arbitrarily chose montmorillonite_1 for this merged file.
The sensitivity of the optical properties to this assumption should be investigated.
The _log10 imaginary index variables reported in EgH79 are omitted.

Reference: EgH79
Egan, W. G., and T. W. Hilgeman (1979), Optical Properties of Inhomogeneous Materials: Applications to Geology, Astronomy, Chemistry, and Engineering, Academic Press, San Diego, CA, 235 pp..

Data from 0.185--2.6 microns measured for illite, kaolinite, montmorillonite
Illite EgH79 p. 103 sample from Fithian, Illinois
Kaolinite EgH79 p. 105 sample from Macon, Georgia
Montmorillonite_I  EgH79 p. 113 sample from Clay Spur, Wyoming
Montmorillonite_II EgH79 p. 115 sample from Amory, Missippippi
Montmorillonite_II has a slightly different wavelength grid than the other minerals
Montmorillonite_II has no measurement at 0.215 um
Montmorillonite_II has a measurement at 0.355 um instead of 0.360 um
These differences are so slight that I placed Montmorillonite_II
on the standard EgH79 wavelength grid by creating an artificial
entry for 0.215 um as the average of the 0.210 and 0.220 entries,
and simply shifting the 0.355 um entry to 0.360 um.

************************************************************************
Begin Procedure to create netCDF from idx_rfr_EgH79 and idx_rfr_roush_* files:
************************************************************************
ncpdq -O --reorder=-bnd -v bnd,idx_rfr_illite_rl,idx_rfr_illite_img -p ${DATA}/aca idx_rfr_roush_illite.nc ~/foo_illite_rdr.nc
ncdump ~/foo_illite_rdr.nc > ~/foo_illite_rdr.cdl
ncpdq -O --reorder=-bnd -v bnd,idx_rfr_kaolinite_rl,idx_rfr_kaolinite_img -p ${DATA}/aca idx_rfr_roush_kaolinite.nc ~/foo_kaolinite_rdr.nc
ncdump ~/foo_kaolinite_rdr.nc > ~/foo_kaolinite_rdr.cdl
ncpdq -O --reorder=-bnd -v bnd,idx_rfr_montmorillonite_rl,idx_rfr_montmorillonite_img -p ${DATA}/aca idx_rfr_roush_montmorillonite.nc ~/foo_montmorillonite_rdr.nc
ncdump ~/foo_montmorillonite_rdr.nc > ~/foo_montmorillonite_rdr.cdl

ncks -v bnd ~/foo_illite_rdr.nc | m
ncks -u -v bnd,idx_rfr_illite_rl,idx_rfr_illite_img -s '%f, ' ~/foo_illite_rdr.nc | m
************************************************************************
End Procedure to create netCDF from idx_rfr_EgH79 and idx_rfr_roush_* files:
************************************************************************
	";

// Begin contents of file:

	float bnd_illite(bnd_illite) ;
		bnd_illite:units = "microns" ;
		bnd_illite:longname = "Band center wavelength, Illite" ;
		bnd_illite:C_format = "%.5g" ;

	float idx_rfr_illite_rl(bnd_illite) ;
		idx_rfr_illite_rl:units = "" ;
		idx_rfr_illite_rl:longname = "Illite refractive index, real part " ;
		idx_rfr_illite_rl:C_format = "%.4g" ;

	float idx_rfr_illite_img(bnd_illite) ;
		idx_rfr_illite_img:units = "" ;
		idx_rfr_illite_img:longname = "Illite refractive index, imag part " ;
		idx_rfr_illite_img:C_format = "%.3g" ;

	float bnd_kaolinite(bnd_kaolinite) ;
		bnd_kaolinite:units = "microns" ;
		bnd_kaolinite:longname = "Band center wavelength, Kaolinite" ;
		bnd_kaolinite:C_format = "%.5g" ;

	float idx_rfr_kaolinite_rl(bnd_kaolinite) ;
		idx_rfr_kaolinite_rl:units = "" ;
		idx_rfr_kaolinite_rl:longname = "Kaolinite refractive index, real part " ;
		idx_rfr_kaolinite_rl:C_format = "%.4g" ;

	float idx_rfr_kaolinite_img(bnd_kaolinite) ;
		idx_rfr_kaolinite_img:units = "" ;
		idx_rfr_kaolinite_img:longname = "Kaolinite refractive index, imag part " ;
		idx_rfr_kaolinite_img:C_format = "%.3g" ;

	float bnd_montmorillonite(bnd_montmorillonite) ;
		bnd_montmorillonite:units = "microns" ;
		bnd_montmorillonite:longname = "Band center wavelength, Montmorillonite" ;
		bnd_montmorillonite:C_format = "%.5g" ;

	float idx_rfr_montmorillonite_rl(bnd_montmorillonite) ;
		idx_rfr_montmorillonite_rl:units = "" ;
		idx_rfr_montmorillonite_rl:longname = "Montmorillonite refractive index, real part " ;
		idx_rfr_montmorillonite_rl:C_format = "%.4g" ;

	float idx_rfr_montmorillonite_img(bnd_montmorillonite) ;
		idx_rfr_montmorillonite_img:units = "" ;
		idx_rfr_montmorillonite_img:longname = "Montmorillonite refractive index, imag part " ;
		idx_rfr_montmorillonite_img:C_format = "%.3g" ;

// End contents EgH79.txt file:

data:

 bnd_illite = 0.185, 0.19, 0.2, 0.21, 0.215, 0.22, 0.225, 0.233, 0.24, 0.26, 0.28, 
    0.3, 0.325, 0.36, 0.37, 0.4, 0.433, 0.466, 0.5, 0.533, 0.566, 0.6, 0.633, 
    0.666, 0.7, 0.817, 0.907, 1, 1.105, 1.2, 1.303, 1.4, 1.5, 1.6, 1.7, 1.8, 
    1.9, 2, 2.1, 2.2, 2.3, 2.4, 2.4999, 
// NB: Relabel EgH79 value at 2.5 um as 2.4999 um to make room for 2.5 um Roush datum
// NB: Excise EgH79 value at 2.6 um in favor of Roush data
// end EgH79 Illite. Begin Roush Illite:
    2.5, 2.5006, 2.5013, 2.5019, 2.5025, 2.5031, 2.5038, 2.5044, 2.505, 
    2.5056, 2.5063, 2.5069, 2.5075, 2.5082, 2.5088, 2.5094, 2.51, 2.5107, 
    2.5113, 2.5119, 2.5126, 2.5132, 2.5138, 2.5145, 2.5151, 2.5157, 2.5164, 
    2.517, 2.5176, 2.5183, 2.5189, 2.5195, 2.5202, 2.5208, 2.5214, 2.5221, 
    2.5227, 2.5233, 2.524, 2.5246, 2.5253, 2.5259, 2.5265, 2.5272, 2.5278, 
    2.5284, 2.5291, 2.5297, 2.5304, 2.531, 2.5316, 2.5323, 2.5329, 2.5336, 
    2.5342, 2.5349, 2.5355, 2.5361, 2.5368, 2.5374, 2.5381, 2.5387, 2.5394, 
    2.54, 2.5407, 2.5413, 2.5419, 2.5426, 2.5432, 2.5439, 2.5445, 2.5452, 
    2.5458, 2.5465, 2.5471, 2.5478, 2.5484, 2.5491, 2.5497, 2.5504, 2.551, 
    2.5517, 2.5523, 2.553, 2.5536, 2.5543, 2.5549, 2.5556, 2.5562, 2.5569, 
    2.5575, 2.5582, 2.5589, 2.5595, 2.5602, 2.5608, 2.5615, 2.5621, 2.5628, 
    2.5634, 2.5641, 2.5648, 2.5654, 2.5661, 2.5667, 2.5674, 2.5681, 2.5687, 
    2.5694, 2.57, 2.5707, 2.5714, 2.572, 2.5727, 2.5733, 2.574, 2.5747, 
    2.5753, 2.576, 2.5767, 2.5773, 2.578, 2.5786, 2.5793, 2.58, 2.5806, 
    2.5813, 2.582, 2.5826, 2.5833, 2.584, 2.5846, 2.5853, 2.586, 2.5867, 
    2.5873, 2.588, 2.5887, 2.5893, 2.59, 2.5907, 2.5913, 2.592, 2.5927, 
    2.5934, 2.594, 2.5947, 2.5954, 2.5961, 2.5967, 2.5974, 2.5981, 2.5988, 
    2.5994, 2.6001, 2.6008, 2.6015, 2.6021, 2.6028, 2.6035, 2.6042, 2.6048, 
    2.6055, 2.6062, 2.6069, 2.6076, 2.6082, 2.6089, 2.6096, 2.6103, 2.611, 
    2.6116, 2.6123, 2.613, 2.6137, 2.6144, 2.6151, 2.6157, 2.6164, 2.6171, 
    2.6178, 2.6185, 2.6192, 2.6199, 2.6205, 2.6212, 2.6219, 2.6226, 2.6233, 
    2.624, 2.6247, 2.6254, 2.6261, 2.6267, 2.6274, 2.6281, 2.6288, 2.6295, 
    2.6302, 2.6309, 2.6316, 2.6323, 2.633, 2.6337, 2.6344, 2.635, 2.6357, 
    2.6364, 2.6371, 2.6378, 2.6385, 2.6392, 2.6399, 2.6406, 2.6413, 2.642, 
    2.6427, 2.6434, 2.6441, 2.6448, 2.6455, 2.6462, 2.6469, 2.6476, 2.6483, 
    2.649, 2.6497, 2.6504, 2.6511, 2.6518, 2.6525, 2.6532, 2.6539, 2.6546, 
    2.6553, 2.656, 2.6567, 2.6575, 2.6582, 2.6589, 2.6596, 2.6603, 2.661, 
    2.6617, 2.6624, 2.6631, 2.6638, 2.6645, 2.6652, 2.666, 2.6667, 2.6674, 
    2.6681, 2.6688, 2.6695, 2.6702, 2.6709, 2.6717, 2.6724, 2.6731, 2.6738, 
    2.6745, 2.6752, 2.6759, 2.6767, 2.6774, 2.6781, 2.6788, 2.6795, 2.6802, 
    2.681, 2.6817, 2.6824, 2.6831, 2.6838, 2.6846, 2.6853, 2.686, 2.6867, 
    2.6874, 2.6882, 2.6889, 2.6896, 2.6903, 2.6911, 2.6918, 2.6925, 2.6932, 
    2.694, 2.6947, 2.6954, 2.6961, 2.6969, 2.6976, 2.6983, 2.6991, 2.6998, 
    2.7005, 2.7012, 2.702, 2.7027, 2.7034, 2.7042, 2.7049, 2.7056, 2.7064, 
    2.7071, 2.7078, 2.7086, 2.7093, 2.71, 2.7108, 2.7115, 2.7122, 2.713, 
    2.7137, 2.7144, 2.7152, 2.7159, 2.7167, 2.7174, 2.7181, 2.7189, 2.7196, 
    2.7203, 2.7211, 2.7218, 2.7226, 2.7233, 2.7241, 2.7248, 2.7255, 2.7263, 
    2.727, 2.7278, 2.7285, 2.7293, 2.73, 2.7307, 2.7315, 2.7322, 2.733, 
    2.7337, 2.7345, 2.7352, 2.736, 2.7367, 2.7375, 2.7382, 2.739, 2.7397, 
    2.7405, 2.7412, 2.742, 2.7427, 2.7435, 2.7442, 2.745, 2.7457, 2.7465, 
    2.7473, 2.748, 2.7488, 2.7495, 2.7503, 2.751, 2.7518, 2.7525, 2.7533, 
    2.7541, 2.7548, 2.7556, 2.7563, 2.7571, 2.7579, 2.7586, 2.7594, 2.7601, 
    2.7609, 2.7617, 2.7624, 2.7632, 2.764, 2.7647, 2.7655, 2.7663, 2.767, 
    2.7678, 2.7685, 2.7693, 2.7701, 2.7709, 2.7716, 2.7724, 2.7732, 2.7739, 
    2.7747, 2.7755, 2.7762, 2.777, 2.7778, 2.7785, 2.7793, 2.7801, 2.7809, 
    2.7816, 2.7824, 2.7832, 2.784, 2.7847, 2.7855, 2.7863, 2.7871, 2.7878, 
    2.7886, 2.7894, 2.7902, 2.791, 2.7917, 2.7925, 2.7933, 2.7941, 2.7949, 
    2.7956, 2.7964, 2.7972, 2.798, 2.7988, 2.7996, 2.8003, 2.8011, 2.8019, 
    2.8027, 2.8035, 2.8043, 2.805, 2.8058, 2.8066, 2.8074, 2.8082, 2.809, 
    2.8098, 2.8106, 2.8114, 2.8121, 2.8129, 2.8137, 2.8145, 2.8153, 2.8161, 
    2.8169, 2.8177, 2.8185, 2.8193, 2.8201, 2.8209, 2.8217, 2.8225, 2.8233, 
    2.8241, 2.8249, 2.8257, 2.8265, 2.8273, 2.8281, 2.8289, 2.8297, 2.8305, 
    2.8313, 2.8321, 2.8329, 2.8337, 2.8345, 2.8353, 2.8361, 2.8369, 2.8377, 
    2.8385, 2.8393, 2.8401, 2.8409, 2.8417, 2.8425, 2.8433, 2.8441, 2.845, 
    2.8458, 2.8466, 2.8474, 2.8482, 2.849, 2.8498, 2.8506, 2.8514, 2.8523, 
    2.8531, 2.8539, 2.8547, 2.8555, 2.8563, 2.8571, 2.858, 2.8588, 2.8596, 
    2.8604, 2.8612, 2.862, 2.8629, 2.8637, 2.8645, 2.8653, 2.8662, 2.867, 
    2.8678, 2.8686, 2.8694, 2.8703, 2.8711, 2.8719, 2.8727, 2.8736, 2.8744, 
    2.8752, 2.876, 2.8769, 2.8777, 2.8785, 2.8794, 2.8802, 2.881, 2.8818, 
    2.8827, 2.8835, 2.8843, 2.8852, 2.886, 2.8868, 2.8877, 2.8885, 2.8893, 
    2.8902, 2.891, 2.8918, 2.8927, 2.8935, 2.8944, 2.8952, 2.896, 2.8969, 
    2.8977, 2.8986, 2.8994, 2.9002, 2.9011, 2.9019, 2.9028, 2.9036, 2.9044, 
    2.9053, 2.9061, 2.907, 2.9078, 2.9087, 2.9095, 2.9104, 2.9112, 2.9121, 
    2.9129, 2.9138, 2.9146, 2.9155, 2.9163, 2.9172, 2.918, 2.9189, 2.9197, 
    2.9206, 2.9214, 2.9223, 2.9231, 2.924, 2.9248, 2.9257, 2.9265, 2.9274, 
    2.9283, 2.9291, 2.93, 2.9308, 2.9317, 2.9326, 2.9334, 2.9343, 2.9351, 
    2.936, 2.9369, 2.9377, 2.9386, 2.9394, 2.9403, 2.9412, 2.942, 2.9429, 
    2.9438, 2.9446, 2.9455, 2.9464, 2.9472, 2.9481, 2.949, 2.9499, 2.9507, 
    2.9516, 2.9525, 2.9533, 2.9542, 2.9551, 2.956, 2.9568, 2.9577, 2.9586, 
    2.9595, 2.9603, 2.9612, 2.9621, 2.963, 2.9638, 2.9647, 2.9656, 2.9665, 
    2.9674, 2.9682, 2.9691, 2.97, 2.9709, 2.9718, 2.9727, 2.9735, 2.9744, 
    2.9753, 2.9762, 2.9771, 2.978, 2.9789, 2.9797, 2.9806, 2.9815, 2.9824, 
    2.9833, 2.9842, 2.9851, 2.986, 2.9869, 2.9878, 2.9886, 2.9895, 2.9904, 
    2.9913, 2.9922, 2.9931, 2.994, 2.9949, 2.9958, 2.9967, 2.9976, 2.9985, 
    2.9994, 3.0003, 3.0012, 3.0021, 3.003, 3.0039, 3.0048, 3.0057, 3.0066, 
    3.0075, 3.0084, 3.0093, 3.0102, 3.0111, 3.012, 3.013, 3.0139, 3.0148, 
    3.0157, 3.0166, 3.0175, 3.0184, 3.0193, 3.0202, 3.0211, 3.0221, 3.023, 
    3.0239, 3.0248, 3.0257, 3.0266, 3.0276, 3.0285, 3.0294, 3.0303, 3.0312, 
    3.0321, 3.0331, 3.034, 3.0349, 3.0358, 3.0367, 3.0377, 3.0386, 3.0395, 
    3.0404, 3.0414, 3.0423, 3.0432, 3.0441, 3.0451, 3.046, 3.0469, 3.0479, 
    3.0488, 3.0497, 3.0506, 3.0516, 3.0525, 3.0534, 3.0544, 3.0553, 3.0562, 
    3.0572, 3.0581, 3.059, 3.06, 3.0609, 3.0618, 3.0628, 3.0637, 3.0647, 
    3.0656, 3.0665, 3.0675, 3.0684, 3.0694, 3.0703, 3.0713, 3.0722, 3.0731, 
    3.0741, 3.075, 3.076, 3.0769, 3.0779, 3.0788, 3.0798, 3.0807, 3.0817, 
    3.0826, 3.0836, 3.0845, 3.0855, 3.0864, 3.0874, 3.0883, 3.0893, 3.0902, 
    3.0912, 3.0921, 3.0931, 3.0941, 3.095, 3.096, 3.0969, 3.0979, 3.0989, 
    3.0998, 3.1008, 3.1017, 3.1027, 3.1037, 3.1046, 3.1056, 3.1066, 3.1075, 
    3.1085, 3.1095, 3.1104, 3.1114, 3.1124, 3.1133, 3.1143, 3.1153, 3.1162, 
    3.1172, 3.1182, 3.1192, 3.1201, 3.1211, 3.1221, 3.123, 3.124, 3.125, 
    3.126, 3.127, 3.1279, 3.1289, 3.1299, 3.1309, 3.1319, 3.1328, 3.1338, 
    3.1348, 3.1358, 3.1368, 3.1377, 3.1387, 3.1397, 3.1407, 3.1417, 3.1427, 
    3.1437, 3.1447, 3.1456, 3.1466, 3.1476, 3.1486, 3.1496, 3.1506, 3.1516, 
    3.1526, 3.1536, 3.1546, 3.1556, 3.1566, 3.1576, 3.1586, 3.1596, 3.1606, 
    3.1616, 3.1626, 3.1636, 3.1646, 3.1656, 3.1666, 3.1676, 3.1686, 3.1696, 
    3.1706, 3.1716, 3.1726, 3.1736, 3.1746, 3.1756, 3.1766, 3.1776, 3.1786, 
    3.1797, 3.1807, 3.1817, 3.1827, 3.1837, 3.1847, 3.1857, 3.1867, 3.1878, 
    3.1888, 3.1898, 3.1908, 3.1918, 3.1928, 3.1939, 3.1949, 3.1959, 3.1969, 
    3.198, 3.199, 3.2, 3.201, 3.202, 3.2031, 3.2041, 3.2051, 3.2062, 3.2072, 
    3.2082, 3.2092, 3.2103, 3.2113, 3.2123, 3.2134, 3.2144, 3.2154, 3.2165, 
    3.2175, 3.2185, 3.2196, 3.2206, 3.2216, 3.2227, 3.2237, 3.2248, 3.2258, 
    3.2268, 3.2279, 3.2289, 3.23, 3.231, 3.2321, 3.2331, 3.2342, 3.2352, 
    3.2362, 3.2373, 3.2383, 3.2394, 3.2404, 3.2415, 3.2425, 3.2436, 3.2446, 
    3.2457, 3.2468, 3.2478, 3.2489, 3.2499, 3.251, 3.252, 3.2531, 3.2541, 
    3.2552, 3.2563, 3.2573, 3.2584, 3.2595, 3.2605, 3.2616, 3.2626, 3.2637, 
    3.2648, 3.2658, 3.2669, 3.268, 3.269, 3.2701, 3.2712, 3.2723, 3.2733, 
    3.2744, 3.2755, 3.2765, 3.2776, 3.2787, 3.2798, 3.2808, 3.2819, 3.283, 
    3.2841, 3.2852, 3.2862, 3.2873, 3.2884, 3.2895, 3.2906, 3.2916, 3.2927, 
    3.2938, 3.2949, 3.296, 3.2971, 3.2982, 3.2992, 3.3003, 3.3014, 3.3025, 
    3.3036, 3.3047, 3.3058, 3.3069, 3.308, 3.3091, 3.3102, 3.3113, 3.3124, 
    3.3135, 3.3146, 3.3156, 3.3167, 3.3179, 3.319, 3.3201, 3.3212, 3.3223, 
    3.3234, 3.3245, 3.3256, 3.3267, 3.3278, 3.3289, 3.33, 3.3311, 3.3322, 
    3.3333, 3.3344, 3.3356, 3.3367, 3.3378, 3.3389, 3.34, 3.3411, 3.3422, 
    3.3434, 3.3445, 3.3456, 3.3467, 3.3478, 3.349, 3.3501, 3.3512, 3.3523, 
    3.3535, 3.3546, 3.3557, 3.3568, 3.358, 3.3591, 3.3602, 3.3613, 3.3625, 
    3.3636, 3.3647, 3.3659, 3.367, 3.3681, 3.3693, 3.3704, 3.3715, 3.3727, 
    3.3738, 3.375, 3.3761, 3.3772, 3.3784, 3.3795, 3.3807, 3.3818, 3.3829, 
    3.3841, 3.3852, 3.3864, 3.3875, 3.3887, 3.3898, 3.391, 3.3921, 3.3933, 
    3.3944, 3.3956, 3.3967, 3.3979, 3.399, 3.4002, 3.4014, 3.4025, 3.4037, 
    3.4048, 3.406, 3.4072, 3.4083, 3.4095, 3.4106, 3.4118, 3.413, 3.4141, 
    3.4153, 3.4165, 3.4176, 3.4188, 3.42, 3.4211, 3.4223, 3.4235, 3.4247, 
    3.4258, 3.427, 3.4282, 3.4294, 3.4305, 3.4317, 3.4329, 3.4341, 3.4352, 
    3.4364, 3.4376, 3.4388, 3.44, 3.4412, 3.4423, 3.4435, 3.4447, 3.4459, 
    3.4471, 3.4483, 3.4495, 3.4507, 3.4518, 3.453, 3.4542, 3.4554, 3.4566, 
    3.4578, 3.459, 3.4602, 3.4614, 3.4626, 3.4638, 3.465, 3.4662, 3.4674, 
    3.4686, 3.4698, 3.471, 3.4722, 3.4734, 3.4746, 3.4758, 3.4771, 3.4783, 
    3.4795, 3.4807, 3.4819, 3.4831, 3.4843, 3.4855, 3.4868, 3.488, 3.4892, 
    3.4904, 3.4916, 3.4928, 3.4941, 3.4953, 3.4965, 3.4977, 3.499, 3.5002, 
    3.5014, 3.5026, 3.5039, 3.5051, 3.5063, 3.5075, 3.5088, 3.51, 3.5112, 
    3.5125, 3.5137, 3.5149, 3.5162, 3.5174, 3.5186, 3.5199, 3.5211, 3.5224, 
    3.5236, 3.5249, 3.5261, 3.5273, 3.5286, 3.5298, 3.5311, 3.5323, 3.5336, 
    3.5348, 3.5361, 3.5373, 3.5386, 3.5398, 3.5411, 3.5423, 3.5436, 3.5448, 
    3.5461, 3.5474, 3.5486, 3.5499, 3.5511, 3.5524, 3.5537, 3.5549, 3.5562, 
    3.5575, 3.5587, 3.56, 3.5613, 3.5625, 3.5638, 3.5651, 3.5663, 3.5676, 
    3.5689, 3.5702, 3.5714, 3.5727, 3.574, 3.5753, 3.5765, 3.5778, 3.5791, 
    3.5804, 3.5817, 3.5829, 3.5842, 3.5855, 3.5868, 3.5881, 3.5894, 3.5907, 
    3.592, 3.5932, 3.5945, 3.5958, 3.5971, 3.5984, 3.5997, 3.601, 3.6023, 
    3.6036, 3.6049, 3.6062, 3.6075, 3.6088, 3.6101, 3.6114, 3.6127, 3.614, 
    3.6153, 3.6166, 3.6179, 3.6193, 3.6206, 3.6219, 3.6232, 3.6245, 3.6258, 
    3.6271, 3.6284, 3.6298, 3.6311, 3.6324, 3.6337, 3.635, 3.6364, 3.6377, 
    3.639, 3.6403, 3.6417, 3.643, 3.6443, 3.6456, 3.647, 3.6483, 3.6496, 
    3.651, 3.6523, 3.6536, 3.655, 3.6563, 3.6576, 3.659, 3.6603, 3.6617, 
    3.663, 3.6643, 3.6657, 3.667, 3.6684, 3.6697, 3.6711, 3.6724, 3.6738, 
    3.6751, 3.6765, 3.6778, 3.6792, 3.6805, 3.6819, 3.6832, 3.6846, 3.686, 
    3.6873, 3.6887, 3.69, 3.6914, 3.6928, 3.6941, 3.6955, 3.6969, 3.6982, 
    3.6996, 3.701, 3.7023, 3.7037, 3.7051, 3.7064, 3.7078, 3.7092, 3.7106, 
    3.712, 3.7133, 3.7147, 3.7161, 3.7175, 3.7189, 3.7202, 3.7216, 3.723, 
    3.7244, 3.7258, 3.7272, 3.7286, 3.73, 3.7313, 3.7327, 3.7341, 3.7355, 
    3.7369, 3.7383, 3.7397, 3.7411, 3.7425, 3.7439, 3.7453, 3.7467, 3.7481, 
    3.7495, 3.7509, 3.7523, 3.7538, 3.7552, 3.7566, 3.758, 3.7594, 3.7608, 
    3.7622, 3.7636, 3.7651, 3.7665, 3.7679, 3.7693, 3.7707, 3.7722, 3.7736, 
    3.775, 3.7764, 3.7779, 3.7793, 3.7807, 3.7821, 3.7836, 3.785, 3.7864, 
    3.7879, 3.7893, 3.7908, 3.7922, 3.7936, 3.7951, 3.7965, 3.7979, 3.7994, 
    3.8008, 3.8023, 3.8037, 3.8052, 3.8066, 3.8081, 3.8095, 3.811, 3.8124, 
    3.8139, 3.8153, 3.8168, 3.8183, 3.8197, 3.8212, 3.8226, 3.8241, 3.8256, 
    3.827, 3.8285, 3.83, 3.8314, 3.8329, 3.8344, 3.8358, 3.8373, 3.8388, 
    3.8402, 3.8417, 3.8432, 3.8447, 3.8462, 3.8476, 3.8491, 3.8506, 3.8521, 
    3.8536, 3.8551, 3.8565, 3.858, 3.8595, 3.861, 3.8625, 3.864, 3.8655, 
    3.867, 3.8685, 3.87, 3.8715, 3.873, 3.8745, 3.876, 3.8775, 3.879, 3.8805, 
    3.882, 3.8835, 3.885, 3.8865, 3.888, 3.8895, 3.8911, 3.8926, 3.8941, 
    3.8956, 3.8971, 3.8986, 3.9002, 3.9017, 3.9032, 3.9047, 3.9063, 3.9078, 
    3.9093, 3.9108, 3.9124, 3.9139, 3.9154, 3.917, 3.9185, 3.92, 3.9216, 
    3.9231, 3.9246, 3.9262, 3.9277, 3.9293, 3.9308, 3.9324, 3.9339, 3.9355, 
    3.937, 3.9386, 3.9401, 3.9417, 3.9432, 3.9448, 3.9463, 3.9479, 3.9494, 
    3.951, 3.9526, 3.9541, 3.9557, 3.9573, 3.9588, 3.9604, 3.962, 3.9635, 
    3.9651, 3.9667, 3.9683, 3.9698, 3.9714, 3.973, 3.9746, 3.9761, 3.9777, 
    3.9793, 3.9809, 3.9825, 3.9841, 3.9857, 3.9872, 3.9888, 3.9904, 3.992, 
    3.9936, 3.9952, 3.9968, 3.9984, 4, 4.0016, 4.0032, 4.0048, 4.0064, 4.008, 
    4.0096, 4.0112, 4.0128, 4.0145, 4.0161, 4.0177, 4.0193, 4.0209, 4.0225, 
    4.0241, 4.0258, 4.0274, 4.029, 4.0306, 4.0323, 4.0339, 4.0355, 4.0371, 
    4.0388, 4.0404, 4.042, 4.0437, 4.0453, 4.0469, 4.0486, 4.0502, 4.0519, 
    4.0535, 4.0552, 4.0568, 4.0584, 4.0601, 4.0617, 4.0634, 4.065, 4.0667, 
    4.0683, 4.07, 4.0717, 4.0733, 4.075, 4.0766, 4.0783, 4.08, 4.0816, 
    4.0833, 4.085, 4.0866, 4.0883, 4.09, 4.0917, 4.0933, 4.095, 4.0967, 
    4.0984, 4.1, 4.1017, 4.1034, 4.1051, 4.1068, 4.1085, 4.1102, 4.1118, 
    4.1135, 4.1152, 4.1169, 4.1186, 4.1203, 4.122, 4.1237, 4.1254, 4.1271, 
    4.1288, 4.1305, 4.1322, 4.1339, 4.1356, 4.1374, 4.1391, 4.1408, 4.1425, 
    4.1442, 4.1459, 4.1477, 4.1494, 4.1511, 4.1528, 4.1545, 4.1563, 4.158, 
    4.1597, 4.1615, 4.1632, 4.1649, 4.1667, 4.1684, 4.1701, 4.1719, 4.1736, 
    4.1754, 4.1771, 4.1789, 4.1806, 4.1824, 4.1841, 4.1859, 4.1876, 4.1894, 
    4.1911, 4.1929, 4.1946, 4.1964, 4.1982, 4.1999, 4.2017, 4.2034, 4.2052, 
    4.207, 4.2088, 4.2105, 4.2123, 4.2141, 4.2159, 4.2176, 4.2194, 4.2212, 
    4.223, 4.2248, 4.2265, 4.2283, 4.2301, 4.2319, 4.2337, 4.2355, 4.2373, 
    4.2391, 4.2409, 4.2427, 4.2445, 4.2463, 4.2481, 4.2499, 4.2517, 4.2535, 
    4.2553, 4.2571, 4.2589, 4.2608, 4.2626, 4.2644, 4.2662, 4.268, 4.2699, 
    4.2717, 4.2735, 4.2753, 4.2772, 4.279, 4.2808, 4.2827, 4.2845, 4.2863, 
    4.2882, 4.29, 4.2918, 4.2937, 4.2955, 4.2974, 4.2992, 4.3011, 4.3029, 
    4.3048, 4.3066, 4.3085, 4.3103, 4.3122, 4.3141, 4.3159, 4.3178, 4.3197, 
    4.3215, 4.3234, 4.3253, 4.3271, 4.329, 4.3309, 4.3328, 4.3346, 4.3365, 
    4.3384, 4.3403, 4.3422, 4.344, 4.3459, 4.3478, 4.3497, 4.3516, 4.3535, 
    4.3554, 4.3573, 4.3592, 4.3611, 4.363, 4.3649, 4.3668, 4.3687, 4.3706, 
    4.3725, 4.3745, 4.3764, 4.3783, 4.3802, 4.3821, 4.384, 4.386, 4.3879, 
    4.3898, 4.3917, 4.3937, 4.3956, 4.3975, 4.3995, 4.4014, 4.4033, 4.4053, 
    4.4072, 4.4092, 4.4111, 4.4131, 4.415, 4.417, 4.4189, 4.4209, 4.4228, 
    4.4248, 4.4267, 4.4287, 4.4307, 4.4326, 4.4346, 4.4366, 4.4385, 4.4405, 
    4.4425, 4.4444, 4.4464, 4.4484, 4.4504, 4.4524, 4.4543, 4.4563, 4.4583, 
    4.4603, 4.4623, 4.4643, 4.4663, 4.4683, 4.4703, 4.4723, 4.4743, 4.4763, 
    4.4783, 4.4803, 4.4823, 4.4843, 4.4863, 4.4883, 4.4903, 4.4924, 4.4944, 
    4.4964, 4.4984, 4.5005, 4.5025, 4.5045, 4.5065, 4.5086, 4.5106, 4.5126, 
    4.5147, 4.5167, 4.5188, 4.5208, 4.5228, 4.5249, 4.5269, 4.529, 4.531, 
    4.5331, 4.5351, 4.5372, 4.5393, 4.5413, 4.5434, 4.5455, 4.5475, 4.5496, 
    4.5517, 4.5537, 4.5558, 4.5579, 4.56, 4.562, 4.5641, 4.5662, 4.5683, 
    4.5704, 4.5725, 4.5746, 4.5767, 4.5788, 4.5809, 4.583, 4.5851, 4.5872, 
    4.5893, 4.5914, 4.5935, 4.5956, 4.5977, 4.5998, 4.6019, 4.6041, 4.6062, 
    4.6083, 4.6104, 4.6125, 4.6147, 4.6168, 4.6189, 4.6211, 4.6232, 4.6253, 
    4.6275, 4.6296, 4.6318, 4.6339, 4.6361, 4.6382, 4.6404, 4.6425, 4.6447, 
    4.6468, 4.649, 4.6512, 4.6533, 4.6555, 4.6577, 4.6598, 4.662, 4.6642, 
    4.6664, 4.6685, 4.6707, 4.6729, 4.6751, 4.6773, 4.6795, 4.6816, 4.6838, 
    4.686, 4.6882, 4.6904, 4.6926, 4.6948, 4.697, 4.6992, 4.7015, 4.7037, 
    4.7059, 4.7081, 4.7103, 4.7125, 4.7148, 4.717, 4.7192, 4.7214, 4.7237, 
    4.7259, 4.7281, 4.7304, 4.7326, 4.7348, 4.7371, 4.7393, 4.7416, 4.7438, 
    4.7461, 4.7483, 4.7506, 4.7529, 4.7551, 4.7574, 4.7596, 4.7619, 4.7642, 
    4.7664, 4.7687, 4.771, 4.7733, 4.7755, 4.7778, 4.7801, 4.7824, 4.7847, 
    4.787, 4.7893, 4.7916, 4.7939, 4.7962, 4.7985, 4.8008, 4.8031, 4.8054, 
    4.8077, 4.81, 4.8123, 4.8146, 4.817, 4.8193, 4.8216, 4.8239, 4.8263, 
    4.8286, 4.8309, 4.8333, 4.8356, 4.8379, 4.8403, 4.8426, 4.845, 4.8473, 
    4.8497, 4.852, 4.8544, 4.8567, 4.8591, 4.8614, 4.8638, 4.8662, 4.8685, 
    4.8709, 4.8733, 4.8757, 4.878, 4.8804, 4.8828, 4.8852, 4.8876, 4.89, 
    4.8924, 4.8948, 4.8972, 4.8996, 4.902, 4.9044, 4.9068, 4.9092, 4.9116, 
    4.914, 4.9164, 4.9188, 4.9213, 4.9237, 4.9261, 4.9285, 4.931, 4.9334, 
    4.9358, 4.9383, 4.9407, 4.9432, 4.9456, 4.948, 4.9505, 4.9529, 4.9554, 
    4.9579, 4.9603, 4.9628, 4.9652, 4.9677, 4.9702, 4.9727, 4.9751, 4.9776, 
    4.9801, 4.9826, 4.985, 4.9875, 4.99, 4.9925, 4.995, 4.9975, 5, 5.0025, 
    5.005, 5.0075, 5.01, 5.0125, 5.015, 5.0176, 5.0201, 5.0226, 5.0251, 
    5.0277, 5.0302, 5.0327, 5.0352, 5.0378, 5.0403, 5.0429, 5.0454, 5.048, 
    5.0505, 5.0531, 5.0556, 5.0582, 5.0607, 5.0633, 5.0659, 5.0684, 5.071, 
    5.0736, 5.0761, 5.0787, 5.0813, 5.0839, 5.0865, 5.0891, 5.0916, 5.0942, 
    5.0968, 5.0994, 5.102, 5.1046, 5.1073, 5.1099, 5.1125, 5.1151, 5.1177, 
    5.1203, 5.123, 5.1256, 5.1282, 5.1308, 5.1335, 5.1361, 5.1387, 5.1414, 
    5.144, 5.1467, 5.1493, 5.152, 5.1546, 5.1573, 5.16, 5.1626, 5.1653, 
    5.168, 5.1706, 5.1733, 5.176, 5.1787, 5.1813, 5.184, 5.1867, 5.1894, 
    5.1921, 5.1948, 5.1975, 5.2002, 5.2029, 5.2056, 5.2083, 5.211, 5.2138, 
    5.2165, 5.2192, 5.2219, 5.2247, 5.2274, 5.2301, 5.2329, 5.2356, 5.2383, 
    5.2411, 5.2438, 5.2466, 5.2493, 5.2521, 5.2549, 5.2576, 5.2604, 5.2632, 
    5.2659, 5.2687, 5.2715, 5.2743, 5.277, 5.2798, 5.2826, 5.2854, 5.2882, 
    5.291, 5.2938, 5.2966, 5.2994, 5.3022, 5.305, 5.3079, 5.3107, 5.3135, 
    5.3163, 5.3191, 5.322, 5.3248, 5.3277, 5.3305, 5.3333, 5.3362, 5.339, 
    5.3419, 5.3447, 5.3476, 5.3505, 5.3533, 5.3562, 5.3591, 5.3619, 5.3648, 
    5.3677, 5.3706, 5.3735, 5.3763, 5.3792, 5.3821, 5.385, 5.3879, 5.3908, 
    5.3937, 5.3967, 5.3996, 5.4025, 5.4054, 5.4083, 5.4113, 5.4142, 5.4171, 
    5.4201, 5.423, 5.4259, 5.4289, 5.4318, 5.4348, 5.4377, 5.4407, 5.4437, 
    5.4466, 5.4496, 5.4526, 5.4555, 5.4585, 5.4615, 5.4645, 5.4675, 5.4705, 
    5.4735, 5.4765, 5.4795, 5.4825, 5.4855, 5.4885, 5.4915, 5.4945, 5.4975, 
    5.5006, 5.5036, 5.5066, 5.5096, 5.5127, 5.5157, 5.5188, 5.5218, 5.5249, 
    5.5279, 5.531, 5.534, 5.5371, 5.5402, 5.5432, 5.5463, 5.5494, 5.5525, 
    5.5556, 5.5586, 5.5617, 5.5648, 5.5679, 5.571, 5.5741, 5.5772, 5.5804, 
    5.5835, 5.5866, 5.5897, 5.5928, 5.596, 5.5991, 5.6022, 5.6054, 5.6085, 
    5.6117, 5.6148, 5.618, 5.6211, 5.6243, 5.6275, 5.6306, 5.6338, 5.637, 
    5.6402, 5.6433, 5.6465, 5.6497, 5.6529, 5.6561, 5.6593, 5.6625, 5.6657, 
    5.6689, 5.6721, 5.6754, 5.6786, 5.6818, 5.685, 5.6883, 5.6915, 5.6948, 
    5.698, 5.7013, 5.7045, 5.7078, 5.711, 5.7143, 5.7176, 5.7208, 5.7241, 
    5.7274, 5.7307, 5.7339, 5.7372, 5.7405, 5.7438, 5.7471, 5.7504, 5.7537, 
    5.7571, 5.7604, 5.7637, 5.767, 5.7703, 5.7737, 5.777, 5.7803, 5.7837, 
    5.787, 5.7904, 5.7937, 5.7971, 5.8005, 5.8038, 5.8072, 5.8106, 5.814, 
    5.8173, 5.8207, 5.8241, 5.8275, 5.8309, 5.8343, 5.8377, 5.8411, 5.8445, 
    5.848, 5.8514, 5.8548, 5.8582, 5.8617, 5.8651, 5.8685, 5.872, 5.8754, 
    5.8789, 5.8824, 5.8858, 5.8893, 5.8928, 5.8962, 5.8997, 5.9032, 5.9067, 
    5.9102, 5.9137, 5.9172, 5.9207, 5.9242, 5.9277, 5.9312, 5.9347, 5.9382, 
    5.9418, 5.9453, 5.9488, 5.9524, 5.9559, 5.9595, 5.963, 5.9666, 5.9701, 
    5.9737, 5.9773, 5.9809, 5.9844, 5.988, 5.9916, 5.9952, 5.9988, 6.0024, 
    6.006, 6.0096, 6.0132, 6.0168, 6.0205, 6.0241, 6.0277, 6.0314, 6.035, 
    6.0386, 6.0423, 6.0459, 6.0496, 6.0533, 6.0569, 6.0606, 6.0643, 6.068, 
    6.0716, 6.0753, 6.079, 6.0827, 6.0864, 6.0901, 6.0938, 6.0976, 6.1013, 
    6.105, 6.1087, 6.1125, 6.1162, 6.12, 6.1237, 6.1275, 6.1312, 6.135, 
    6.1387, 6.1425, 6.1463, 6.1501, 6.1538, 6.1576, 6.1614, 6.1652, 6.169, 
    6.1728, 6.1767, 6.1805, 6.1843, 6.1881, 6.192, 6.1958, 6.1996, 6.2035, 
    6.2073, 6.2112, 6.215, 6.2189, 6.2228, 6.2267, 6.2305, 6.2344, 6.2383, 
    6.2422, 6.2461, 6.25, 6.2539, 6.2578, 6.2617, 6.2657, 6.2696, 6.2735, 
    6.2775, 6.2814, 6.2854, 6.2893, 6.2933, 6.2972, 6.3012, 6.3052, 6.3091, 
    6.3131, 6.3171, 6.3211, 6.3251, 6.3291, 6.3331, 6.3371, 6.3412, 6.3452, 
    6.3492, 6.3532, 6.3573, 6.3613, 6.3654, 6.3694, 6.3735, 6.3776, 6.3816, 
    6.3857, 6.3898, 6.3939, 6.398, 6.402, 6.4061, 6.4103, 6.4144, 6.4185, 
    6.4226, 6.4267, 6.4309, 6.435, 6.4392, 6.4433, 6.4475, 6.4516, 6.4558, 
    6.4599, 6.4641, 6.4683, 6.4725, 6.4767, 6.4809, 6.4851, 6.4893, 6.4935, 
    6.4977, 6.502, 6.5062, 6.5104, 6.5147, 6.5189, 6.5232, 6.5274, 6.5317, 
    6.5359, 6.5402, 6.5445, 6.5488, 6.5531, 6.5574, 6.5617, 6.566, 6.5703, 
    6.5746, 6.5789, 6.5833, 6.5876, 6.592, 6.5963, 6.6007, 6.605, 6.6094, 
    6.6138, 6.6181, 6.6225, 6.6269, 6.6313, 6.6357, 6.6401, 6.6445, 6.6489, 
    6.6534, 6.6578, 6.6622, 6.6667, 6.6711, 6.6756, 6.68, 6.6845, 6.689, 
    6.6934, 6.6979, 6.7024, 6.7069, 6.7114, 6.7159, 6.7204, 6.7249, 6.7295, 
    6.734, 6.7385, 6.7431, 6.7476, 6.7522, 6.7568, 6.7613, 6.7659, 6.7705, 
    6.7751, 6.7797, 6.7843, 6.7889, 6.7935, 6.7981, 6.8027, 6.8074, 6.812, 
    6.8166, 6.8213, 6.8259, 6.8306, 6.8353, 6.8399, 6.8446, 6.8493, 6.854, 
    6.8587, 6.8634, 6.8681, 6.8729, 6.8776, 6.8823, 6.8871, 6.8918, 6.8966, 
    6.9013, 6.9061, 6.9109, 6.9156, 6.9204, 6.9252, 6.93, 6.9348, 6.9396, 
    6.9444, 6.9493, 6.9541, 6.9589, 6.9638, 6.9686, 6.9735, 6.9784, 6.9832, 
    6.9881, 6.993, 6.9979, 7.0028, 7.0077, 7.0126, 7.0175, 7.0225, 7.0274, 
    7.0323, 7.0373, 7.0423, 7.0472, 7.0522, 7.0572, 7.0621, 7.0671, 7.0721, 
    7.0771, 7.0822, 7.0872, 7.0922, 7.0972, 7.1023, 7.1073, 7.1124, 7.1174, 
    7.1225, 7.1276, 7.1327, 7.1378, 7.1429, 7.148, 7.1531, 7.1582, 7.1633, 
    7.1685, 7.1736, 7.1788, 7.1839, 7.1891, 7.1942, 7.1994, 7.2046, 7.2098, 
    7.215, 7.2202, 7.2254, 7.2307, 7.2359, 7.2411, 7.2464, 7.2516, 7.2569, 
    7.2622, 7.2674, 7.2727, 7.278, 7.2833, 7.2886, 7.2939, 7.2993, 7.3046, 
    7.3099, 7.3153, 7.3206, 7.326, 7.3314, 7.3368, 7.3421, 7.3475, 7.3529, 
    7.3584, 7.3638, 7.3692, 7.3746, 7.3801, 7.3855, 7.391, 7.3964, 7.4019, 
    7.4074, 7.4129, 7.4184, 7.4239, 7.4294, 7.4349, 7.4405, 7.446, 7.4516, 
    7.4571, 7.4627, 7.4683, 7.4738, 7.4794, 7.485, 7.4906, 7.4963, 7.5019, 
    7.5075, 7.5131, 7.5188, 7.5245, 7.5301, 7.5358, 7.5415, 7.5472, 7.5529, 
    7.5586, 7.5643, 7.57, 7.5758, 7.5815, 7.5873, 7.593, 7.5988, 7.6046, 
    7.6104, 7.6161, 7.622, 7.6278, 7.6336, 7.6394, 7.6453, 7.6511, 7.657, 
    7.6628, 7.6687, 7.6746, 7.6805, 7.6864, 7.6923, 7.6982, 7.7042, 7.7101, 
    7.716, 7.722, 7.728, 7.734, 7.7399, 7.7459, 7.7519, 7.758, 7.764, 7.77, 
    7.776, 7.7821, 7.7882, 7.7942, 7.8003, 7.8064, 7.8125, 7.8186, 7.8247, 
    7.8309, 7.837, 7.8431, 7.8493, 7.8555, 7.8616, 7.8678, 7.874, 7.8802, 
    7.8864, 7.8927, 7.8989, 7.9051, 7.9114, 7.9177, 7.9239, 7.9302, 7.9365, 
    7.9428, 7.9491, 7.9554, 7.9618, 7.9681, 7.9745, 7.9808, 7.9872, 7.9936, 
    8, 8.0064, 8.0128, 8.0192, 8.0257, 8.0321, 8.0386, 8.0451, 8.0515, 8.058, 
    8.0645, 8.071, 8.0775, 8.0841, 8.0906, 8.0972, 8.1037, 8.1103, 8.1169, 
    8.1235, 8.1301, 8.1367, 8.1433, 8.15, 8.1566, 8.1633, 8.1699, 8.1766, 
    8.1833, 8.19, 8.1967, 8.2034, 8.2102, 8.2169, 8.2237, 8.2305, 8.2372, 
    8.244, 8.2508, 8.2576, 8.2645, 8.2713, 8.2781, 8.285, 8.2919, 8.2988, 
    8.3056, 8.3126, 8.3195, 8.3264, 8.3333, 8.3403, 8.3472, 8.3542, 8.3612, 
    8.3682, 8.3752, 8.3822, 8.3893, 8.3963, 8.4034, 8.4104, 8.4175, 8.4246, 
    8.4317, 8.4388, 8.4459, 8.4531, 8.4602, 8.4674, 8.4746, 8.4818, 8.489, 
    8.4962, 8.5034, 8.5106, 8.5179, 8.5251, 8.5324, 8.5397, 8.547, 8.5543, 
    8.5616, 8.569, 8.5763, 8.5837, 8.5911, 8.5985, 8.6059, 8.6133, 8.6207, 
    8.6281, 8.6356, 8.643, 8.6505, 8.658, 8.6655, 8.673, 8.6806, 8.6881, 
    8.6957, 8.7032, 8.7108, 8.7184, 8.726, 8.7336, 8.7413, 8.7489, 8.7566, 
    8.7642, 8.7719, 8.7796, 8.7873, 8.7951, 8.8028, 8.8106, 8.8183, 8.8261, 
    8.8339, 8.8417, 8.8496, 8.8574, 8.8652, 8.8731, 8.881, 8.8889, 8.8968, 
    8.9047, 8.9127, 8.9206, 8.9286, 8.9366, 8.9445, 8.9526, 8.9606, 8.9686, 
    8.9767, 8.9847, 8.9928, 9.0009, 9.009, 9.0171, 9.0253, 9.0334, 9.0416, 
    9.0498, 9.058, 9.0662, 9.0744, 9.0827, 9.0909, 9.0992, 9.1075, 9.1158, 
    9.1241, 9.1324, 9.1408, 9.1491, 9.1575, 9.1659, 9.1743, 9.1827, 9.1912, 
    9.1996, 9.2081, 9.2166, 9.2251, 9.2336, 9.2421, 9.2507, 9.2593, 9.2678, 
    9.2764, 9.2851, 9.2937, 9.3023, 9.311, 9.3197, 9.3284, 9.3371, 9.3458, 
    9.3545, 9.3633, 9.3721, 9.3809, 9.3897, 9.3985, 9.4073, 9.4162, 9.4251, 
    9.434, 9.4429, 9.4518, 9.4607, 9.4697, 9.4787, 9.4877, 9.4967, 9.5057, 
    9.5147, 9.5238, 9.5329, 9.542, 9.5511, 9.5602, 9.5694, 9.5785, 9.5877, 
    9.5969, 9.6061, 9.6154, 9.6246, 9.6339, 9.6432, 9.6525, 9.6618, 9.6712, 
    9.6805, 9.6899, 9.6993, 9.7087, 9.7182, 9.7276, 9.7371, 9.7466, 9.7561, 
    9.7656, 9.7752, 9.7847, 9.7943, 9.8039, 9.8135, 9.8232, 9.8328, 9.8425, 
    9.8522, 9.8619, 9.8717, 9.8814, 9.8912, 9.901, 9.9108, 9.9206, 9.9305, 
    9.9404, 9.9502, 9.9602, 9.9701, 9.98, 9.99, 10, 10.01, 10.02, 10.03, 
    10.04, 10.05, 10.06, 10.071, 10.081, 10.091, 10.101, 10.111, 10.122, 
    10.132, 10.142, 10.152, 10.163, 10.173, 10.183, 10.194, 10.204, 10.215, 
    10.225, 10.235, 10.246, 10.256, 10.267, 10.278, 10.288, 10.299, 10.309, 
    10.32, 10.331, 10.341, 10.352, 10.363, 10.373, 10.384, 10.395, 10.406, 
    10.417, 10.427, 10.438, 10.449, 10.46, 10.471, 10.482, 10.493, 10.504, 
    10.515, 10.526, 10.537, 10.549, 10.56, 10.571, 10.582, 10.593, 10.604, 
    10.616, 10.627, 10.638, 10.65, 10.661, 10.672, 10.684, 10.695, 10.707, 
    10.718, 10.73, 10.741, 10.753, 10.764, 10.776, 10.788, 10.799, 10.811, 
    10.823, 10.834, 10.846, 10.858, 10.87, 10.881, 10.893, 10.905, 10.917, 
    10.929, 10.941, 10.953, 10.965, 10.977, 10.989, 11.001, 11.013, 11.025, 
    11.038, 11.05, 11.062, 11.074, 11.087, 11.099, 11.111, 11.123, 11.136, 
    11.148, 11.161, 11.173, 11.186, 11.198, 11.211, 11.223, 11.236, 11.249, 
    11.261, 11.274, 11.287, 11.299, 11.312, 11.325, 11.338, 11.351, 11.364, 
    11.377, 11.389, 11.403, 11.415, 11.429, 11.442, 11.455, 11.468, 11.481, 
    11.494, 11.507, 11.521, 11.534, 11.547, 11.561, 11.574, 11.587, 11.601, 
    11.614, 11.628, 11.641, 11.655, 11.669, 11.682, 11.696, 11.71, 11.723, 
    11.737, 11.751, 11.765, 11.779, 11.792, 11.806, 11.82, 11.834, 11.848, 
    11.862, 11.877, 11.891, 11.905, 11.919, 11.933, 11.947, 11.962, 11.976, 
    11.99, 12.005, 12.019, 12.034, 12.048, 12.063, 12.077, 12.092, 12.106, 
    12.121, 12.136, 12.151, 12.165, 12.18, 12.195, 12.21, 12.225, 12.24, 
    12.255, 12.27, 12.285, 12.3, 12.315, 12.33, 12.346, 12.361, 12.376, 
    12.392, 12.407, 12.422, 12.438, 12.453, 12.469, 12.484, 12.5, 12.516, 
    12.531, 12.547, 12.563, 12.579, 12.594, 12.61, 12.626, 12.642, 12.658, 
    12.674, 12.69, 12.707, 12.723, 12.739, 12.755, 12.771, 12.788, 12.804, 
    12.821, 12.837, 12.854, 12.87, 12.887, 12.903, 12.92, 12.937, 12.953, 
    12.97, 12.987, 13.004, 13.021, 13.038, 13.055, 13.072, 13.089, 13.106, 
    13.123, 13.141, 13.158, 13.175, 13.193, 13.21, 13.227, 13.245, 13.263, 
    13.28, 13.298, 13.316, 13.333, 13.351, 13.369, 13.387, 13.405, 13.423, 
    13.441, 13.459, 13.477, 13.495, 13.514, 13.532, 13.55, 13.568, 13.587, 
    13.605, 13.624, 13.643, 13.661, 13.68, 13.699, 13.717, 13.736, 13.755, 
    13.774, 13.793, 13.812, 13.831, 13.85, 13.87, 13.889, 13.908, 13.928, 
    13.947, 13.967, 13.986, 14.006, 14.025, 14.045, 14.065, 14.085, 14.104, 
    14.124, 14.144, 14.164, 14.184, 14.205, 14.225, 14.245, 14.265, 14.286, 
    14.306, 14.327, 14.347, 14.368, 14.389, 14.409, 14.43, 14.451, 14.472, 
    14.493, 14.514, 14.535, 14.556, 14.577, 14.599, 14.62, 14.641, 14.663, 
    14.684, 14.706, 14.727, 14.749, 14.771, 14.793, 14.815, 14.837, 14.859, 
    14.881, 14.903, 14.925, 14.948, 14.97, 14.993, 15.015, 15.038, 15.06, 
    15.083, 15.106, 15.129, 15.151, 15.175, 15.198, 15.221, 15.244, 15.267, 
    15.29, 15.314, 15.337, 15.361, 15.385, 15.408, 15.432, 15.456, 15.48, 
    15.504, 15.528, 15.552, 15.576, 15.601, 15.625, 15.649, 15.674, 15.699, 
    15.723, 15.748, 15.773, 15.798, 15.823, 15.848, 15.873, 15.898, 15.924, 
    15.949, 15.974, 16, 16.026, 16.051, 16.077, 16.103, 16.129, 16.155, 
    16.181, 16.208, 16.234, 16.26, 16.287, 16.313, 16.34, 16.367, 16.393, 
    16.42, 16.447, 16.475, 16.502, 16.529, 16.556, 16.584, 16.611, 16.639, 
    16.667, 16.694, 16.722, 16.75, 16.778, 16.807, 16.835, 16.863, 16.892, 
    16.92, 16.949, 16.978, 17.007, 17.036, 17.065, 17.094, 17.123, 17.153, 
    17.182, 17.212, 17.241, 17.271, 17.301, 17.331, 17.361, 17.391, 17.422, 
    17.452, 17.483, 17.513, 17.544, 17.575, 17.606, 17.637, 17.668, 17.699, 
    17.73, 17.762, 17.794, 17.825, 17.857, 17.889, 17.921, 17.953, 17.986, 
    18.018, 18.051, 18.083, 18.116, 18.149, 18.182, 18.215, 18.248, 18.281, 
    18.315, 18.349, 18.382, 18.416, 18.45, 18.484, 18.518, 18.553, 18.587, 
    18.622, 18.657, 18.692, 18.727, 18.762, 18.797, 18.832, 18.868, 18.904, 
    18.939, 18.975, 19.011, 19.048, 19.084, 19.121, 19.157, 19.194, 19.231, 
    19.268, 19.305, 19.342, 19.38, 19.417, 19.455, 19.493, 19.531, 19.569, 
    19.608, 19.646, 19.685, 19.724, 19.763, 19.802, 19.841, 19.881, 19.92, 
    19.96, 20, 20.04, 20.08, 20.121, 20.161, 20.202, 20.243, 20.284, 20.325, 
    20.367, 20.408, 20.45, 20.492, 20.534, 20.576, 20.619, 20.661, 20.704, 
    20.747, 20.79, 20.833, 20.877, 20.92, 20.964, 21.008, 21.053, 21.097, 
    21.142, 21.186, 21.231, 21.277, 21.322, 21.368, 21.413, 21.459, 21.505, 
    21.552, 21.598, 21.645, 21.692, 21.739, 21.787, 21.834, 21.882, 21.93, 
    21.978, 22.026, 22.075, 22.124, 22.173, 22.222, 22.272, 22.321, 22.371, 
    22.421, 22.472, 22.522, 22.573, 22.624, 22.676, 22.727, 22.779, 22.831, 
    22.883, 22.936, 22.989, 23.042, 23.095, 23.148, 23.202, 23.256, 23.31, 
    23.365, 23.419, 23.474, 23.529, 23.585, 23.641, 23.697, 23.753, 23.809, 
    23.866, 23.923, 23.981, 24.038, 24.096, 24.155, 24.213, 24.272, 24.331, 
    24.39, 24.45, 24.51, 24.57, 24.631, 24.691, 24.753, 24.814, 24.876, 
    24.938, 25, 25.063, 25.126, 25.189, 25.253, 25.316, 25.381, 25.445, 
    25.51, 25.575, 25.641, 25.707, 25.773, 25.84, 25.907, 25.974, 26.042, 
    26.11, 26.178, 26.247, 26.316, 26.385, 26.455, 26.525, 26.596, 26.667, 
    26.738, 26.81, 26.882, 26.954, 27.027, 27.1, 27.174, 27.248, 27.322, 
    27.397, 27.472, 27.548, 27.624, 27.701, 27.778, 27.855, 27.933, 28.011, 
    28.09, 28.169, 28.249, 28.329, 28.409, 28.49, 28.571, 28.653, 28.736, 
    28.818, 28.902, 28.986, 29.07, 29.154, 29.24, 29.326, 29.412, 29.499, 
    29.586, 29.674, 29.762, 29.851, 29.94, 30.03, 30.121, 30.212, 30.303, 
    30.395, 30.488, 30.581, 30.675, 30.769, 30.864, 30.96, 31.056, 31.153, 
    31.25, 31.348, 31.447, 31.546, 31.646, 31.746, 31.847, 31.949, 32.051, 
    32.154, 32.258, 32.362, 32.467, 32.573, 32.68, 32.787, 32.895, 33.003, 
    33.113, 33.223, 33.333, 33.445, 33.557, 33.67, 33.784, 33.898, 34.014, 
    34.13, 34.247, 34.364, 34.483, 34.602, 34.722, 34.843, 34.965, 35.088, 
    35.211, 35.336, 35.461, 35.587, 35.714, 35.842, 35.971, 36.101, 36.232, 
    36.364, 36.496, 36.63, 36.765, 36.9, 37.037, 37.175, 37.313, 37.453, 
    37.594, 37.736, 37.879, 38.023, 38.168, 38.314, 38.461, 38.61, 38.76, 
    38.91, 39.062, 39.216, 39.37, 39.526, 39.682, 39.841, 40, 40.161, 40.323, 
    40.486, 40.65, 40.816, 40.984, 41.152, 41.322, 41.494, 41.667, 41.841, 
    42.017, 42.194, 42.373, 42.553, 42.735, 42.918, 43.103, 43.29, 43.478, 
    43.668, 43.86, 44.053, 44.248, 44.444, 44.643, 44.843, 45.045, 45.249, 
    45.454, 45.662, 45.872, 46.083, 46.296, 46.512, 46.729, 46.948, 47.17, 
    47.393, 47.619, 47.847, 48.077, 48.309, 48.544, 48.78, 49.02, 49.261, 
    49.505, 49.751, 50, 50.251, 50.505, 50.761, 51.02, 51.282, 51.546, 
    51.813, 52.083, 52.356, 52.632, 52.91, 53.192, 53.476, 53.763, 54.054, 
    54.348, 54.645, 54.945, 55.249, 55.556, 55.866, 56.18, 56.497, 56.818, 
    57.143, 57.471, 57.804, 58.139, 58.479, 58.824, 59.172, 59.524, 59.88, 
    60.241, 60.606, 60.976, 61.35, 61.728, 62.112, 62.5, 62.893, 63.291, 
    63.694, 64.103, 64.516, 64.935, 65.359, 65.789, 66.225, 66.667, 67.114, 
    67.568, 68.027, 68.493, 68.965, 69.444, 69.93, 70.423, 70.922, 71.429, 
    71.942, 72.464, 72.993, 73.529, 74.074, 74.627, 75.188, 75.758, 76.336, 
    76.923, 77.519, 78.125, 78.74, 79.365, 80, 80.645, 81.301, 81.967, 
    82.645, 83.333, 84.034, 84.746, 85.47, 86.207, 86.956, 87.719, 88.496, 
    89.286, 90.09, 90.909, 91.743, 92.593, 93.458, 94.34, 95.238, 96.154, 
    97.087, 98.039, 99.01, 100, 101.01, 102.04, 103.09, 104.17, 105.26, 
    106.38, 107.53, 108.7, 109.89, 111.11, 112.36, 113.64, 114.94, 116.28, 
    117.65, 119.05, 120.48, 121.95, 123.46, 125, 126.58, 128.21, 129.87, 
    131.58, 133.33, 135.14, 136.99, 138.89, 140.85, 142.86, 144.93, 147.06, 
    149.25, 151.52, 153.85, 156.25, 158.73, 161.29, 163.93, 166.67, 169.49, 
    172.41, 175.44, 178.57, 181.82, 185.19, 188.68, 192.31, 196.08, 200 ;

 idx_rfr_illite_rl = 1.448, 1.444, 1.441, 1.438, 1.434, 1.431, 1.427, 1.424, 
    1.42, 1.417, 1.411, 1.401, 1.404, 1.406, 1.415, 1.423, 1.42, 1.418, 
    1.415, 1.414, 1.412, 1.411, 1.407, 1.403, 1.399, 1.395, 1.391, 1.387, 
    1.387, 1.387, 1.387, 1.387, 1.387, 1.387, 1.387, 1.387, 1.387, 1.387, 
    1.387, 1.387, 1.387, 1.387, 1.387,
// NB: Relabel EgH79 value at 2.5 um as 2.4999 um to make room for 2.5 um Roush datum
// NB: Excise EgH79 value at 2.6 um in favor of Roush data
// end EgH79 Illite. Begin Roush Illite:
    1.381, 1.381, 1.381, 1.381, 1.381, 1.381, 1.38, 1.38, 
    1.38, 1.381, 1.381, 1.381, 1.381, 1.381, 1.381, 1.381, 1.382, 1.382, 
    1.382, 1.382, 1.382, 1.382, 1.382, 1.381, 1.381, 1.381, 1.38, 1.38, 1.38, 
    1.38, 1.38, 1.38, 1.38, 1.38, 1.38, 1.38, 1.381, 1.381, 1.382, 1.382, 
    1.383, 1.383, 1.384, 1.384, 1.384, 1.384, 1.384, 1.384, 1.384, 1.385, 
    1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 
    1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 
    1.385, 1.384, 1.384, 1.383, 1.383, 1.382, 1.382, 1.382, 1.382, 1.381, 
    1.381, 1.381, 1.381, 1.381, 1.381, 1.381, 1.382, 1.382, 1.383, 1.384, 
    1.384, 1.385, 1.385, 1.385, 1.384, 1.384, 1.383, 1.382, 1.382, 1.381, 
    1.38, 1.38, 1.38, 1.38, 1.38, 1.38, 1.381, 1.381, 1.381, 1.381, 1.381, 
    1.381, 1.381, 1.381, 1.381, 1.38, 1.38, 1.381, 1.381, 1.381, 1.381, 
    1.382, 1.383, 1.383, 1.384, 1.384, 1.384, 1.384, 1.383, 1.383, 1.382, 
    1.382, 1.381, 1.38, 1.38, 1.38, 1.38, 1.381, 1.381, 1.382, 1.382, 1.383, 
    1.383, 1.383, 1.383, 1.383, 1.382, 1.382, 1.382, 1.381, 1.381, 1.381, 
    1.381, 1.382, 1.382, 1.382, 1.382, 1.382, 1.382, 1.381, 1.38, 1.379, 
    1.378, 1.377, 1.376, 1.375, 1.375, 1.375, 1.376, 1.377, 1.378, 1.379, 
    1.381, 1.382, 1.383, 1.384, 1.384, 1.384, 1.383, 1.382, 1.382, 1.38, 
    1.379, 1.378, 1.378, 1.378, 1.378, 1.378, 1.379, 1.38, 1.381, 1.381, 
    1.382, 1.382, 1.382, 1.382, 1.381, 1.381, 1.38, 1.379, 1.379, 1.378, 
    1.378, 1.377, 1.377, 1.377, 1.377, 1.378, 1.378, 1.378, 1.378, 1.379, 
    1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.379, 1.379, 1.379, 1.378, 1.378, 1.378, 
    1.378, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.378, 
    1.378, 1.378, 1.379, 1.379, 1.38, 1.38, 1.379, 1.379, 1.379, 1.378, 
    1.378, 1.377, 1.376, 1.375, 1.374, 1.373, 1.372, 1.371, 1.37, 1.369, 
    1.369, 1.368, 1.368, 1.367, 1.367, 1.367, 1.367, 1.367, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.367, 1.367, 1.367, 1.366, 
    1.366, 1.365, 1.365, 1.364, 1.363, 1.363, 1.362, 1.361, 1.36, 1.36, 
    1.359, 1.358, 1.358, 1.358, 1.357, 1.357, 1.356, 1.356, 1.356, 1.355, 
    1.355, 1.355, 1.355, 1.354, 1.354, 1.353, 1.353, 1.352, 1.35, 1.349, 
    1.349, 1.348, 1.347, 1.346, 1.346, 1.346, 1.346, 1.346, 1.346, 1.346, 
    1.346, 1.346, 1.345, 1.345, 1.344, 1.343, 1.342, 1.341, 1.34, 1.339, 
    1.339, 1.338, 1.338, 1.338, 1.338, 1.339, 1.34, 1.34, 1.341, 1.342, 
    1.342, 1.343, 1.343, 1.343, 1.343, 1.342, 1.342, 1.341, 1.34, 1.34, 
    1.339, 1.339, 1.338, 1.338, 1.339, 1.339, 1.34, 1.34, 1.342, 1.343, 
    1.344, 1.345, 1.347, 1.348, 1.349, 1.35, 1.351, 1.352, 1.352, 1.352, 
    1.353, 1.353, 1.353, 1.354, 1.355, 1.356, 1.357, 1.358, 1.36, 1.361, 
    1.362, 1.364, 1.365, 1.365, 1.366, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.368, 1.368, 1.368, 1.369, 1.369, 1.37, 1.371, 1.371, 1.372, 1.373, 
    1.374, 1.375, 1.376, 1.376, 1.377, 1.378, 1.378, 1.378, 1.378, 1.379, 
    1.378, 1.378, 1.378, 1.378, 1.377, 1.377, 1.376, 1.376, 1.376, 1.375, 
    1.375, 1.375, 1.374, 1.374, 1.374, 1.373, 1.373, 1.372, 1.372, 1.371, 
    1.371, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.371, 1.371, 1.371, 
    1.372, 1.372, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.374, 
    1.373, 1.373, 1.373, 1.372, 1.372, 1.371, 1.371, 1.37, 1.369, 1.369, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.369, 1.369, 1.369, 1.37, 1.37, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.37, 1.37, 1.37, 1.369, 1.368, 1.368, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.368, 1.368, 1.368, 1.369, 1.369, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.366, 1.366, 
    1.366, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.372, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 
    1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 1.363, 1.363, 1.363, 
    1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 
    1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.362, 1.362, 1.362, 
    1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 
    1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.361, 1.361, 1.361, 
    1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 
    1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.36, 1.36, 1.36, 1.36, 
    1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.359, 
    1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 
    1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.358, 
    1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.357, 
    1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.356, 
    1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 
    1.355, 1.355, 1.355, 1.356, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 
    1.355, 1.355, 1.355, 1.355, 1.354, 1.354, 1.354, 1.354, 1.354, 1.354, 
    1.354, 1.354, 1.354, 1.354, 1.353, 1.353, 1.353, 1.353, 1.353, 1.353, 
    1.353, 1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 
    1.352, 1.351, 1.351, 1.351, 1.351, 1.351, 1.351, 1.351, 1.351, 1.35, 
    1.35, 1.35, 1.35, 1.35, 1.35, 1.35, 1.349, 1.349, 1.349, 1.349, 1.349, 
    1.348, 1.348, 1.348, 1.348, 1.348, 1.348, 1.348, 1.348, 1.348, 1.347, 
    1.347, 1.347, 1.347, 1.347, 1.347, 1.346, 1.346, 1.346, 1.346, 1.346, 
    1.346, 1.346, 1.345, 1.345, 1.345, 1.345, 1.345, 1.345, 1.344, 1.344, 
    1.344, 1.344, 1.344, 1.344, 1.344, 1.344, 1.344, 1.343, 1.343, 1.343, 
    1.343, 1.343, 1.343, 1.342, 1.342, 1.342, 1.342, 1.342, 1.341, 1.341, 
    1.341, 1.341, 1.341, 1.341, 1.341, 1.341, 1.34, 1.34, 1.34, 1.34, 1.34, 
    1.34, 1.34, 1.34, 1.339, 1.339, 1.34, 1.339, 1.339, 1.339, 1.339, 1.339, 
    1.339, 1.339, 1.338, 1.338, 1.338, 1.338, 1.338, 1.338, 1.337, 1.337, 
    1.337, 1.337, 1.337, 1.336, 1.336, 1.336, 1.336, 1.336, 1.336, 1.336, 
    1.335, 1.335, 1.335, 1.335, 1.335, 1.335, 1.334, 1.334, 1.334, 1.334, 
    1.334, 1.334, 1.334, 1.334, 1.334, 1.334, 1.333, 1.333, 1.333, 1.333, 
    1.333, 1.333, 1.333, 1.332, 1.332, 1.332, 1.332, 1.332, 1.332, 1.332, 
    1.332, 1.331, 1.331, 1.331, 1.331, 1.331, 1.331, 1.331, 1.33, 1.33, 1.33, 
    1.33, 1.33, 1.33, 1.33, 1.33, 1.329, 1.329, 1.329, 1.329, 1.329, 1.329, 
    1.329, 1.329, 1.329, 1.328, 1.328, 1.328, 1.328, 1.328, 1.328, 1.327, 
    1.327, 1.327, 1.327, 1.327, 1.327, 1.327, 1.326, 1.326, 1.326, 1.326, 
    1.326, 1.326, 1.326, 1.326, 1.325, 1.325, 1.325, 1.325, 1.325, 1.325, 
    1.325, 1.325, 1.325, 1.325, 1.324, 1.324, 1.324, 1.324, 1.324, 1.324, 
    1.324, 1.324, 1.324, 1.324, 1.324, 1.324, 1.324, 1.323, 1.323, 1.323, 
    1.323, 1.322, 1.322, 1.322, 1.322, 1.322, 1.322, 1.322, 1.322, 1.322, 
    1.322, 1.322, 1.322, 1.321, 1.321, 1.321, 1.321, 1.321, 1.321, 1.321, 
    1.321, 1.32, 1.32, 1.32, 1.32, 1.32, 1.32, 1.32, 1.32, 1.319, 1.319, 
    1.319, 1.319, 1.319, 1.319, 1.319, 1.319, 1.319, 1.319, 1.319, 1.319, 
    1.319, 1.319, 1.319, 1.318, 1.318, 1.318, 1.318, 1.318, 1.318, 1.317, 
    1.317, 1.317, 1.317, 1.317, 1.317, 1.317, 1.317, 1.316, 1.316, 1.316, 
    1.316, 1.316, 1.316, 1.316, 1.316, 1.315, 1.315, 1.315, 1.315, 1.315, 
    1.315, 1.315, 1.315, 1.314, 1.314, 1.314, 1.314, 1.314, 1.314, 1.314, 
    1.313, 1.313, 1.313, 1.313, 1.313, 1.312, 1.312, 1.312, 1.312, 1.312, 
    1.312, 1.312, 1.311, 1.311, 1.311, 1.311, 1.311, 1.311, 1.31, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.309, 1.309, 1.309, 1.309, 1.309, 
    1.309, 1.309, 1.308, 1.308, 1.308, 1.308, 1.308, 1.308, 1.307, 1.307, 
    1.307, 1.307, 1.307, 1.306, 1.306, 1.306, 1.306, 1.306, 1.305, 1.305, 
    1.305, 1.305, 1.305, 1.305, 1.305, 1.305, 1.305, 1.305, 1.304, 1.304, 
    1.304, 1.304, 1.304, 1.304, 1.304, 1.303, 1.303, 1.303, 1.303, 1.303, 
    1.303, 1.302, 1.302, 1.302, 1.302, 1.302, 1.302, 1.301, 1.301, 1.301, 
    1.301, 1.301, 1.301, 1.3, 1.3, 1.3, 1.3, 1.3, 1.299, 1.299, 1.299, 1.299, 
    1.299, 1.298, 1.298, 1.298, 1.298, 1.297, 1.297, 1.297, 1.297, 1.297, 
    1.297, 1.296, 1.296, 1.296, 1.296, 1.296, 1.295, 1.295, 1.295, 1.295, 
    1.295, 1.294, 1.294, 1.294, 1.294, 1.294, 1.294, 1.293, 1.293, 1.293, 
    1.293, 1.293, 1.293, 1.293, 1.292, 1.292, 1.292, 1.292, 1.291, 1.291, 
    1.291, 1.291, 1.29, 1.29, 1.29, 1.29, 1.289, 1.289, 1.289, 1.289, 1.289, 
    1.288, 1.288, 1.288, 1.288, 1.287, 1.287, 1.287, 1.287, 1.286, 1.286, 
    1.286, 1.285, 1.285, 1.285, 1.285, 1.284, 1.284, 1.284, 1.283, 1.283, 
    1.283, 1.282, 1.282, 1.282, 1.282, 1.281, 1.281, 1.281, 1.28, 1.28, 1.28, 
    1.28, 1.279, 1.279, 1.279, 1.279, 1.278, 1.278, 1.278, 1.278, 1.277, 
    1.277, 1.276, 1.276, 1.276, 1.275, 1.275, 1.275, 1.274, 1.274, 1.274, 
    1.273, 1.273, 1.273, 1.273, 1.272, 1.272, 1.271, 1.271, 1.271, 1.27, 
    1.27, 1.27, 1.269, 1.269, 1.269, 1.268, 1.268, 1.268, 1.267, 1.267, 
    1.266, 1.266, 1.266, 1.266, 1.265, 1.265, 1.265, 1.264, 1.264, 1.263, 
    1.263, 1.263, 1.262, 1.262, 1.262, 1.261, 1.261, 1.26, 1.26, 1.26, 1.259, 
    1.259, 1.258, 1.258, 1.258, 1.258, 1.258, 1.257, 1.257, 1.257, 1.256, 
    1.256, 1.256, 1.255, 1.255, 1.255, 1.255, 1.254, 1.254, 1.253, 1.253, 
    1.253, 1.252, 1.252, 1.251, 1.251, 1.251, 1.251, 1.251, 1.25, 1.25, 
    1.249, 1.249, 1.249, 1.249, 1.248, 1.248, 1.247, 1.247, 1.247, 1.247, 
    1.246, 1.246, 1.246, 1.245, 1.245, 1.245, 1.245, 1.244, 1.244, 1.244, 
    1.244, 1.244, 1.244, 1.243, 1.243, 1.242, 1.242, 1.242, 1.242, 1.241, 
    1.241, 1.24, 1.24, 1.24, 1.24, 1.239, 1.239, 1.239, 1.238, 1.238, 1.238, 
    1.237, 1.237, 1.237, 1.237, 1.237, 1.237, 1.236, 1.236, 1.236, 1.235, 
    1.235, 1.235, 1.235, 1.234, 1.235, 1.234, 1.234, 1.233, 1.233, 1.233, 
    1.233, 1.232, 1.232, 1.231, 1.231, 1.231, 1.231, 1.23, 1.23, 1.23, 1.229, 
    1.229, 1.229, 1.228, 1.228, 1.228, 1.228, 1.227, 1.227, 1.226, 1.226, 
    1.226, 1.226, 1.225, 1.225, 1.225, 1.224, 1.224, 1.223, 1.223, 1.222, 
    1.222, 1.222, 1.221, 1.221, 1.221, 1.22, 1.22, 1.219, 1.219, 1.218, 
    1.218, 1.218, 1.217, 1.217, 1.216, 1.215, 1.215, 1.214, 1.214, 1.213, 
    1.213, 1.212, 1.212, 1.211, 1.211, 1.211, 1.21, 1.209, 1.209, 1.208, 
    1.208, 1.207, 1.207, 1.206, 1.205, 1.205, 1.204, 1.204, 1.203, 1.202, 
    1.201, 1.201, 1.2, 1.199, 1.198, 1.198, 1.197, 1.196, 1.195, 1.194, 
    1.194, 1.193, 1.192, 1.191, 1.19, 1.189, 1.188, 1.187, 1.186, 1.185, 
    1.185, 1.183, 1.183, 1.181, 1.181, 1.179, 1.179, 1.177, 1.177, 1.175, 
    1.174, 1.173, 1.171, 1.171, 1.169, 1.168, 1.167, 1.166, 1.165, 1.165, 
    1.164, 1.163, 1.162, 1.162, 1.16, 1.159, 1.158, 1.157, 1.156, 1.154, 
    1.153, 1.151, 1.15, 1.148, 1.147, 1.146, 1.145, 1.144, 1.143, 1.142, 
    1.141, 1.14, 1.139, 1.138, 1.136, 1.135, 1.135, 1.134, 1.133, 1.132, 
    1.131, 1.13, 1.129, 1.127, 1.126, 1.125, 1.122, 1.12, 1.118, 1.116, 
    1.114, 1.112, 1.11, 1.109, 1.107, 1.106, 1.105, 1.104, 1.104, 1.102, 
    1.101, 1.101, 1.099, 1.097, 1.095, 1.093, 1.091, 1.089, 1.086, 1.084, 
    1.082, 1.079, 1.077, 1.075, 1.072, 1.071, 1.068, 1.066, 1.063, 1.06, 
    1.057, 1.053, 1.051, 1.048, 1.045, 1.042, 1.04, 1.038, 1.036, 1.035, 
    1.033, 1.032, 1.03, 1.03, 1.028, 1.027, 1.025, 1.023, 1.02, 1.017, 1.014, 
    1.01, 1.008, 1.004, 1, 0.997, 0.994, 0.99, 0.987, 0.984, 0.981, 0.978, 
    0.974, 0.971, 0.968, 0.964, 0.96, 0.957, 0.952, 0.948, 0.944, 0.94, 
    0.936, 0.932, 0.928, 0.925, 0.921, 0.917, 0.914, 0.91, 0.907, 0.903, 0.9, 
    0.897, 0.893, 0.889, 0.886, 0.882, 0.878, 0.874, 0.871, 0.867, 0.864, 
    0.861, 0.858, 0.855, 0.852, 0.849, 0.846, 0.843, 0.84, 0.837, 0.834, 
    0.831, 0.827, 0.824, 0.82, 0.816, 0.812, 0.808, 0.805, 0.801, 0.797, 
    0.793, 0.788, 0.784, 0.78, 0.776, 0.772, 0.768, 0.764, 0.76, 0.756, 
    0.752, 0.749, 0.747, 0.744, 0.743, 0.742, 0.742, 0.743, 0.744, 0.745, 
    0.746, 0.747, 0.747, 0.747, 0.745, 0.742, 0.739, 0.734, 0.729, 0.723, 
    0.716, 0.71, 0.703, 0.698, 0.692, 0.688, 0.684, 0.681, 0.679, 0.678, 
    0.677, 0.676, 0.676, 0.677, 0.677, 0.678, 0.679, 0.68, 0.682, 0.683, 
    0.685, 0.686, 0.688, 0.69, 0.691, 0.693, 0.695, 0.697, 0.7, 0.702, 0.704, 
    0.706, 0.708, 0.71, 0.712, 0.715, 0.717, 0.719, 0.722, 0.724, 0.727, 
    0.729, 0.732, 0.735, 0.738, 0.741, 0.744, 0.748, 0.751, 0.755, 0.76, 
    0.764, 0.769, 0.774, 0.779, 0.785, 0.79, 0.797, 0.803, 0.81, 0.817, 
    0.824, 0.831, 0.839, 0.846, 0.853, 0.861, 0.868, 0.875, 0.882, 0.889, 
    0.896, 0.902, 0.908, 0.914, 0.919, 0.924, 0.93, 0.935, 0.94, 0.945, 0.95, 
    0.955, 0.96, 0.965, 0.971, 0.976, 0.982, 0.987, 0.993, 0.999, 1.005, 
    1.011, 1.017, 1.023, 1.03, 1.037, 1.045, 1.053, 1.062, 1.072, 1.083, 
    1.095, 1.108, 1.122, 1.137, 1.154, 1.172, 1.192, 1.213, 1.236, 1.26, 
    1.285, 1.312, 1.34, 1.37, 1.4, 1.431, 1.463, 1.495, 1.528, 1.56, 1.592, 
    1.623, 1.653, 1.683, 1.711, 1.738, 1.764, 1.789, 1.812, 1.835, 1.856, 
    1.876, 1.895, 1.913, 1.931, 1.948, 1.965, 1.981, 1.997, 2.012, 2.028, 
    2.042, 2.057, 2.072, 2.086, 2.101, 2.115, 2.128, 2.142, 2.155, 2.168, 
    2.181, 2.192, 2.204, 2.214, 2.224, 2.233, 2.242, 2.249, 2.256, 2.262, 
    2.268, 2.273, 2.277, 2.281, 2.285, 2.288, 2.29, 2.292, 2.293, 2.294, 
    2.294, 2.292, 2.291, 2.288, 2.284, 2.279, 2.273, 2.266, 2.258, 2.25, 
    2.241, 2.231, 2.22, 2.209, 2.198, 2.187, 2.175, 2.163, 2.151, 2.139, 
    2.126, 2.114, 2.101, 2.089, 2.076, 2.064, 2.052, 2.039, 2.027, 2.015, 
    2.003, 1.991, 1.98, 1.969, 1.958, 1.947, 1.937, 1.927, 1.917, 1.908, 
    1.899, 1.891, 1.883, 1.876, 1.868, 1.862, 1.855, 1.849, 1.843, 1.838, 
    1.833, 1.828, 1.824, 1.82, 1.817, 1.814, 1.811, 1.809, 1.807, 1.805, 
    1.804, 1.803, 1.803, 1.803, 1.803, 1.804, 1.805, 1.807, 1.808, 1.811, 
    1.813, 1.815, 1.818, 1.82, 1.822, 1.824, 1.825, 1.826, 1.825, 1.825, 
    1.823, 1.821, 1.818, 1.814, 1.809, 1.805, 1.799, 1.794, 1.788, 1.782, 
    1.776, 1.771, 1.766, 1.761, 1.756, 1.751, 1.747, 1.743, 1.739, 1.736, 
    1.732, 1.729, 1.725, 1.721, 1.718, 1.714, 1.71, 1.706, 1.703, 1.699, 
    1.695, 1.692, 1.688, 1.684, 1.681, 1.677, 1.674, 1.67, 1.666, 1.663, 
    1.659, 1.655, 1.651, 1.648, 1.644, 1.641, 1.637, 1.633, 1.63, 1.626, 
    1.623, 1.619, 1.616, 1.612, 1.608, 1.605, 1.601, 1.597, 1.593, 1.589, 
    1.586, 1.582, 1.579, 1.576, 1.573, 1.571, 1.568, 1.566, 1.565, 1.563, 
    1.562, 1.56, 1.558, 1.557, 1.555, 1.553, 1.551, 1.548, 1.546, 1.543, 
    1.539, 1.535, 1.531, 1.527, 1.521, 1.515, 1.509, 1.502, 1.494, 1.485, 
    1.477, 1.468, 1.46, 1.451, 1.444, 1.438, 1.434, 1.431, 1.43, 1.431, 
    1.433, 1.438, 1.444, 1.451, 1.458, 1.466, 1.473, 1.479, 1.484, 1.488, 
    1.489, 1.489, 1.488, 1.485, 1.482, 1.479, 1.476, 1.474, 1.474, 1.474, 
    1.476, 1.479, 1.483, 1.489, 1.494, 1.5, 1.505, 1.51, 1.514, 1.517, 1.519, 
    1.519, 1.519, 1.517, 1.515, 1.512, 1.509, 1.506, 1.503, 1.501, 1.499, 
    1.496, 1.495, 1.493, 1.493, 1.492, 1.491, 1.491, 1.491, 1.492, 1.492, 
    1.492, 1.493, 1.493, 1.493, 1.493, 1.492, 1.492, 1.491, 1.489, 1.487, 
    1.485, 1.483, 1.48, 1.478, 1.475, 1.472, 1.469, 1.466, 1.463, 1.461, 
    1.458, 1.456, 1.454, 1.452, 1.45, 1.448, 1.446, 1.444, 1.442, 1.439, 
    1.437, 1.434, 1.431, 1.428, 1.425, 1.422, 1.418, 1.415, 1.412, 1.409, 
    1.405, 1.401, 1.398, 1.394, 1.391, 1.387, 1.383, 1.379, 1.376, 1.372, 
    1.369, 1.366, 1.365, 1.364, 1.363, 1.363, 1.364, 1.365, 1.367, 1.369, 
    1.37, 1.372, 1.372, 1.373, 1.373, 1.373, 1.372, 1.371, 1.369, 1.367, 
    1.364, 1.362, 1.36, 1.357, 1.355, 1.353, 1.35, 1.348, 1.345, 1.343, 
    1.341, 1.338, 1.335, 1.332, 1.329, 1.325, 1.322, 1.318, 1.314, 1.311, 
    1.306, 1.302, 1.298, 1.294, 1.289, 1.285, 1.281, 1.277, 1.273, 1.269, 
    1.265, 1.261, 1.257, 1.253, 1.249, 1.245, 1.242, 1.238, 1.234, 1.23, 
    1.227, 1.223, 1.219, 1.215, 1.212, 1.208, 1.204, 1.201, 1.197, 1.194, 
    1.19, 1.188, 1.184, 1.181, 1.178, 1.175, 1.171, 1.168, 1.163, 1.159, 
    1.154, 1.149, 1.143, 1.137, 1.131, 1.125, 1.119, 1.112, 1.106, 1.1, 
    1.093, 1.087, 1.08, 1.074, 1.067, 1.06, 1.054, 1.047, 1.04, 1.034, 1.027, 
    1.021, 1.014, 1.008, 1.001, 0.995, 0.989, 0.983, 0.978, 0.972, 0.967, 
    0.962, 0.957, 0.953, 0.949, 0.945, 0.941, 0.938, 0.935, 0.933, 0.93, 
    0.928, 0.927, 0.925, 0.924, 0.923, 0.923, 0.922, 0.922, 0.922, 0.923, 
    0.923, 0.924, 0.925, 0.927, 0.929, 0.931, 0.933, 0.936, 0.939, 0.942, 
    0.946, 0.95, 0.954, 0.959, 0.963, 0.968, 0.973, 0.979, 0.984, 0.991, 
    0.997, 1.004, 1.012, 1.021, 1.03, 1.041, 1.052, 1.065, 1.078, 1.093, 
    1.109, 1.125, 1.143, 1.162, 1.181, 1.201, 1.221, 1.242, 1.263, 1.284, 
    1.305, 1.326, 1.346, 1.366, 1.386, 1.404, 1.422, 1.44, 1.456, 1.471, 
    1.486, 1.499, 1.51, 1.521, 1.53, 1.537, 1.542, 1.545, 1.547, 1.546, 
    1.544, 1.54, 1.535, 1.529, 1.521, 1.513, 1.504, 1.496, 1.486, 1.477, 
    1.469, 1.46, 1.452, 1.445, 1.438, 1.432, 1.428, 1.425, 1.423, 1.422, 
    1.424, 1.428, 1.434, 1.443, 1.454, 1.469, 1.486, 1.508, 1.533, 1.561, 
    1.594, 1.63, 1.67, 1.714, 1.76, 1.81, 1.861, 1.913, 1.967, 2.019, 2.07, 
    2.119, 2.164, 2.205, 2.242, 2.274, 2.3, 2.322, 2.34, 2.354, 2.364, 2.372, 
    2.378, 2.382, 2.385, 2.388, 2.391, 2.392, 2.393, 2.394, 2.393, 2.39, 
    2.387, 2.381, 2.374, 2.366, 2.357, 2.347, 2.337, 2.328, 2.319, 2.31, 
    2.303, 2.298, 2.295, 2.293, 2.294, 2.296, 2.3, 2.306, 2.313, 2.322, 
    2.331, 2.341, 2.352, 2.363, 2.373, 2.383, 2.392, 2.401, 2.408, 2.414, 
    2.418, 2.422, 2.423, 2.423, 2.421, 2.417, 2.411, 2.402, 2.39, 2.376, 
    2.36, 2.342, 2.324, 2.306, 2.289, 2.273, 2.261, 2.252, 2.246, 2.245, 
    2.248, 2.253, 2.262, 2.271, 2.282, 2.291, 2.298, 2.301, 2.302, 2.298, 
    2.29, 2.278, 2.264, 2.248, 2.231, 2.214, 2.197, 2.182, 2.17, 2.159, 
    2.152, 2.147, 2.145, 2.146, 2.15, 2.156, 2.164, 2.174, 2.185, 2.196, 
    2.207, 2.217, 2.227, 2.234, 2.24, 2.245, 2.249, 2.252, 2.254, 2.256, 
    2.258, 2.261, 2.264, 2.267, 2.271, 2.276, 2.28, 2.284, 2.288, 2.291, 
    2.294, 2.296, 2.296, 2.296, 2.295, 2.292, 2.289, 2.284, 2.28, 2.274, 
    2.269, 2.263, 2.257, 2.252, 2.247, 2.242, 2.237, 2.233, 2.23, 2.226, 
    2.223, 2.219, 2.216, 2.213, 2.21, 2.207, 2.204, 2.201, 2.199, 2.197, 
    2.195, 2.192, 2.19, 2.188, 2.185, 2.182, 2.18, 2.177, 2.174, 2.171, 
    2.168, 2.164, 2.161, 2.158, 2.154, 2.15, 2.147, 2.143, 2.138, 2.134, 
    2.13, 2.126, 2.122, 2.118, 2.114, 2.11, 2.106, 2.102, 2.099, 2.096, 
    2.092, 2.088, 2.085, 2.081, 2.078, 2.074, 2.07, 2.066, 2.062, 2.058, 
    2.054, 2.049, 2.044, 2.04, 2.036, 2.032, 2.03, 2.028, 2.026, 2.027, 
    2.028, 2.03, 2.034, 2.039, 2.044, 2.051, 2.057, 2.065, 2.072, 2.079, 
    2.086, 2.093, 2.1, 2.106, 2.112, 2.117, 2.122, 2.126, 2.129, 2.132, 
    2.134, 2.136, 2.136, 2.136, 2.135, 2.134, 2.131, 2.128, 2.124, 2.12, 
    2.115, 2.111, 2.107, 2.104, 2.101, 2.097, 2.094, 2.091, 2.088, 2.085, 
    2.081, 2.077, 2.074, 2.072, 2.07, 2.067, 2.065, 2.063, 2.06, 2.057, 
    2.053, 2.05, 2.047, 2.045, 2.044, 2.042, 2.041, 2.039, 2.036, 2.034, 
    2.031, 2.027, 2.023, 2.019, 2.015, 2.012, 2.009, 2.006, 2.003, 2.001, 
    1.999, 1.999, 1.999, 1.999, 2, 2.001, 2.002, 2.004, 2.006, 2.009, 2.012, 
    2.015, 2.02, 2.024, 2.029, 2.033, 2.037, 2.039, 2.041, 2.041, 2.041, 
    2.04, 2.039, 2.037, 2.034, 2.032, 2.029, 2.025, 2.022, 2.018, 2.014, 
    2.01, 2.006, 2.003, 2, 1.997, 1.996, 1.995, 1.994, 1.995, 1.995, 1.995, 
    1.995, 1.995, 1.994, 1.993, 1.992, 1.99, 1.988, 1.986, 1.985, 1.983, 
    1.982, 1.98, 1.979, 1.978, 1.976, 1.975, 1.974, 1.972, 1.972, 1.971, 
    1.971, 1.973, 1.975, 1.978, 1.982, 1.986, 1.99, 1.993, 1.997, 1.999, 
    2.001, 2.002, 2.003, 2.003, 2.002, 2.003, 2.002, 2.002, 2.001, 2, 1.998, 
    1.996, 1.995, 1.996, 1.999, 2.005, 2.015, 2.028, 2.043, 2.06, 2.078, 
    2.097, 2.114, 2.13, 2.145, 2.159, 2.174, 2.187, 2.201, 2.214, 2.227, 
    2.24, 2.254, 2.268, 2.28, 2.291, 2.303, 2.313, 2.322, 2.331, 2.338, 
    2.343, 2.348, 2.353, 2.356, 2.357, 2.355, 2.352, 2.346, 2.339, 2.33, 
    2.322, 2.312, 2.303, 2.296, 2.289, 2.282, 2.274, 2.267, 2.259, 2.252, 
    2.245, 2.239, 2.233, 2.228, 2.224, 2.221, 2.217, 2.214, 2.21, 2.206, 
    2.202, 2.199, 2.196, 2.194, 2.191, 2.19, 2.188 ;

 idx_rfr_illite_img = 0.002238721, 0.002187761, 0.002290867, 0.002344228, 
    0.002398834, 0.002691535, 0.002398834, 0.002344228, 0.002454709, 
    0.002041738, 0.001862087, 0.001819701, 0.001659587, 0.00144544, 
    0.001230269, 0.001174897, 0.001071519, 0.001071519, 0.001023293, 
    0.0008317639, 0.0007079456, 0.0007079456, 0.0006918308, 0.001148153, 
    0.001202264, 0.001230269, 0.001202264, 0.001230269, 0.001174897, 
    0.001174897, 0.001202264, 0.001174897, 0.001148153, 0.001288249, 
    0.001698244, 0.00144544, 0.001778279, 0.001288249, 0.001584893, 
    0.001949844, 0.002691535, 0.002041738, 0.003467368, 
// NB: Relabel EgH79 value at 2.5 um as 2.4999 um to make room for 2.5 um Roush datum
// NB: Excise EgH79 value at 2.6 um in favor of Roush data
// end EgH79 Illite. Begin Roush Illite:
    0.004, 0.004, 0.004, 0.004, 0.005, 0.004, 0.005, 0.005, 
    0.005, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 
    0.006, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.006, 0.006, 
    0.006, 0.007, 0.007, 0.007, 0.008, 0.008, 0.008, 0.009, 0.009, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.009, 0.009, 0.009, 0.009, 0.009, 0.008, 0.008, 
    0.008, 0.008, 0.008, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 
    0.007, 0.007, 0.006, 0.006, 0.006, 0.006, 0.005, 0.005, 0.005, 0.004, 
    0.004, 0.004, 0.003, 0.003, 0.003, 0.003, 0.003, 0.004, 0.004, 0.004, 
    0.004, 0.005, 0.005, 0.006, 0.006, 0.007, 0.007, 0.007, 0.008, 0.008, 
    0.007, 0.007, 0.006, 0.005, 0.005, 0.004, 0.004, 0.003, 0.003, 0.003, 
    0.003, 0.004, 0.004, 0.005, 0.005, 0.006, 0.006, 0.006, 0.006, 0.006, 
    0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.007, 0.007, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.007, 0.006, 0.006, 0.005, 0.005, 
    0.004, 0.004, 0.004, 0.004, 0.005, 0.006, 0.006, 0.006, 0.007, 0.007, 
    0.007, 0.007, 0.007, 0.006, 0.006, 0.005, 0.005, 0.004, 0.004, 0.004, 
    0.004, 0.005, 0.005, 0.005, 0.005, 0.005, 0.004, 0.004, 0.003, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.003, 0.004, 0.006, 0.007, 0.008, 
    0.009, 0.01, 0.01, 0.01, 0.01, 0.009, 0.007, 0.006, 0.005, 0.004, 0.003, 
    0.002, 0.002, 0.003, 0.003, 0.004, 0.005, 0.005, 0.006, 0.007, 0.006, 
    0.006, 0.006, 0.005, 0.005, 0.004, 0.003, 0.003, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.003, 0.003, 0.004, 0.004, 0.005, 0.005, 0.005, 
    0.005, 0.005, 0.004, 0.004, 0.004, 0.004, 0.004, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.002, 0.002, 0.002, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.001, 0.001, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001, 0.002, 0.003, 0.004, 0.005, 
    0.005, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.007, 0.008, 
    0.009, 0.01, 0.011, 0.013, 0.014, 0.016, 0.017, 0.019, 0.02, 0.021, 
    0.021, 0.021, 0.022, 0.022, 0.022, 0.021, 0.021, 0.022, 0.022, 0.022, 
    0.023, 0.024, 0.025, 0.027, 0.028, 0.03, 0.031, 0.033, 0.034, 0.036, 
    0.037, 0.038, 0.039, 0.04, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.042, 0.043, 0.043, 0.044, 0.045, 0.045, 0.046, 
    0.046, 0.046, 0.046, 0.045, 0.044, 0.044, 0.043, 0.043, 0.042, 0.042, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.04, 0.04, 0.039, 0.039, 0.038, 0.037, 0.036, 0.035, 
    0.034, 0.033, 0.032, 0.031, 0.03, 0.03, 0.029, 0.028, 0.028, 0.028, 
    0.027, 0.027, 0.027, 0.027, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 
    0.026, 0.026, 0.026, 0.026, 0.026, 0.027, 0.027, 0.028, 0.028, 0.029, 
    0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.028, 0.028, 0.027, 0.027, 
    0.027, 0.026, 0.026, 0.025, 0.025, 0.024, 0.024, 0.024, 0.023, 0.023, 
    0.023, 0.024, 0.024, 0.025, 0.025, 0.026, 0.026, 0.027, 0.027, 0.028, 
    0.028, 0.028, 0.028, 0.027, 0.027, 0.027, 0.026, 0.025, 0.025, 0.025, 
    0.024, 0.024, 0.025, 0.025, 0.025, 0.026, 0.026, 0.027, 0.027, 0.028, 
    0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.027, 0.027, 0.027, 0.027, 
    0.027, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.027, 0.026, 
    0.026, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 
    0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.028, 0.028, 
    0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 
    0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 
    0.028, 0.028, 0.028, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 
    0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 
    0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.033, 0.033, 0.033, 0.033, 
    0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 
    0.033, 0.033, 0.033, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 
    0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.035, 0.035, 0.035, 
    0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 
    0.035, 0.035, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 
    0.036, 0.036, 0.037, 0.036, 0.036, 0.036, 0.036, 0.037, 0.037, 0.037, 
    0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 
    0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.04, 0.04, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.044, 0.044, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.045, 0.045, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.049, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.05, 0.05, 0.05, 
    0.049, 0.049, 0.049, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.05, 0.05, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.047, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.048, 0.048, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.046, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.045, 0.044, 0.044, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.043, 0.044, 0.044, 0.044, 
    0.043, 0.043, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.043, 0.043, 0.044, 0.044, 0.044, 0.043, 0.043, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.043, 0.043, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.044, 
    0.044, 0.044, 0.044, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.042, 0.043, 0.043, 0.043, 0.042, 0.042, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.042, 0.042, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.041, 0.042, 0.042, 0.042, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.04, 0.04, 0.041, 0.041, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.039, 0.04, 0.04, 0.04, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.038, 0.038, 0.039, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.039, 0.039, 0.039, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.039, 0.039, 0.039, 0.039, 0.038, 
    0.039, 0.039, 0.038, 0.038, 0.039, 0.038, 0.038, 0.039, 0.038, 0.038, 
    0.038, 0.038, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.04, 0.04, 0.039, 
    0.039, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.041, 0.04, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.044, 0.044, 0.043, 0.043, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.046, 0.045, 0.045, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.048, 0.048, 0.048, 0.047, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.049, 0.048, 
    0.048, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.05, 0.049, 0.049, 0.05, 0.05, 
    0.05, 0.049, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.051, 0.051, 
    0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 
    0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 
    0.051, 0.051, 0.051, 0.051, 0.052, 0.051, 0.051, 0.052, 0.051, 0.051, 
    0.052, 0.052, 0.051, 0.052, 0.052, 0.051, 0.052, 0.052, 0.052, 0.052, 
    0.052, 0.052, 0.052, 0.052, 0.052, 0.053, 0.053, 0.053, 0.053, 0.052, 
    0.053, 0.053, 0.052, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.055, 0.055, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.056, 0.055, 0.056, 0.056, 
    0.056, 0.056, 0.055, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 
    0.056, 0.056, 0.056, 0.056, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 
    0.057, 0.057, 0.057, 0.057, 0.057, 0.058, 0.058, 0.058, 0.058, 0.058, 
    0.058, 0.058, 0.058, 0.058, 0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 
    0.059, 0.059, 0.059, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.061, 0.061, 
    0.061, 0.061, 0.062, 0.062, 0.062, 0.062, 0.062, 0.062, 0.062, 0.063, 
    0.063, 0.063, 0.063, 0.063, 0.063, 0.063, 0.063, 0.064, 0.064, 0.064, 
    0.064, 0.064, 0.065, 0.065, 0.065, 0.065, 0.065, 0.065, 0.066, 0.066, 
    0.066, 0.066, 0.066, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.068, 
    0.068, 0.068, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.07, 
    0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.071, 0.071, 0.071, 
    0.071, 0.071, 0.071, 0.071, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 
    0.073, 0.073, 0.073, 0.073, 0.073, 0.074, 0.073, 0.074, 0.074, 0.074, 
    0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 
    0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.075, 0.074, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 
    0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 
    0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 
    0.073, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.071, 
    0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.07, 0.07, 0.07, 0.07, 0.07, 
    0.069, 0.069, 0.069, 0.069, 0.069, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.066, 
    0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 
    0.066, 0.066, 0.066, 0.067, 0.067, 0.067, 0.067, 0.067, 0.068, 0.068, 
    0.068, 0.067, 0.067, 0.067, 0.067, 0.067, 0.066, 0.066, 0.066, 0.066, 
    0.067, 0.067, 0.067, 0.068, 0.068, 0.068, 0.069, 0.069, 0.069, 0.069, 
    0.069, 0.069, 0.069, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.069, 0.069, 
    0.068, 0.068, 0.067, 0.066, 0.066, 0.066, 0.066, 0.067, 0.067, 0.068, 
    0.069, 0.07, 0.071, 0.071, 0.072, 0.071, 0.071, 0.071, 0.071, 0.069, 
    0.069, 0.068, 0.068, 0.067, 0.067, 0.067, 0.068, 0.067, 0.067, 0.068, 
    0.067, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.069, 0.071, 
    0.071, 0.073, 0.074, 0.076, 0.078, 0.08, 0.081, 0.082, 0.083, 0.083, 
    0.085, 0.084, 0.084, 0.084, 0.083, 0.082, 0.083, 0.082, 0.082, 0.083, 
    0.083, 0.084, 0.085, 0.086, 0.086, 0.088, 0.088, 0.09, 0.091, 0.092, 
    0.093, 0.094, 0.094, 0.096, 0.097, 0.098, 0.1, 0.102, 0.104, 0.106, 
    0.108, 0.111, 0.113, 0.116, 0.118, 0.121, 0.123, 0.126, 0.129, 0.132, 
    0.134, 0.137, 0.139, 0.142, 0.145, 0.148, 0.152, 0.155, 0.159, 0.162, 
    0.166, 0.17, 0.173, 0.177, 0.18, 0.184, 0.187, 0.19, 0.194, 0.197, 0.2, 
    0.203, 0.206, 0.21, 0.214, 0.217, 0.221, 0.225, 0.229, 0.234, 0.238, 
    0.243, 0.248, 0.253, 0.258, 0.264, 0.269, 0.275, 0.282, 0.289, 0.296, 
    0.303, 0.311, 0.319, 0.327, 0.335, 0.343, 0.35, 0.356, 0.361, 0.366, 
    0.37, 0.373, 0.375, 0.377, 0.379, 0.381, 0.384, 0.388, 0.392, 0.398, 
    0.404, 0.412, 0.421, 0.431, 0.441, 0.452, 0.462, 0.473, 0.484, 0.495, 
    0.506, 0.516, 0.527, 0.537, 0.546, 0.556, 0.565, 0.575, 0.584, 0.593, 
    0.602, 0.611, 0.62, 0.628, 0.637, 0.646, 0.654, 0.663, 0.671, 0.679, 
    0.688, 0.696, 0.704, 0.713, 0.721, 0.73, 0.738, 0.747, 0.756, 0.764, 
    0.773, 0.782, 0.791, 0.8, 0.81, 0.819, 0.829, 0.838, 0.848, 0.857, 0.867, 
    0.877, 0.886, 0.896, 0.906, 0.915, 0.924, 0.934, 0.942, 0.951, 0.959, 
    0.968, 0.975, 0.983, 0.99, 0.997, 1, 1.01, 1.02, 1.02, 1.03, 1.03, 1.04, 
    1.04, 1.05, 1.06, 1.06, 1.07, 1.08, 1.09, 1.09, 1.1, 1.11, 1.12, 1.12, 
    1.13, 1.14, 1.15, 1.16, 1.17, 1.18, 1.19, 1.2, 1.21, 1.23, 1.24, 1.25, 
    1.27, 1.28, 1.3, 1.31, 1.33, 1.34, 1.36, 1.38, 1.39, 1.41, 1.42, 1.44, 
    1.46, 1.47, 1.48, 1.49, 1.5, 1.51, 1.52, 1.53, 1.53, 1.53, 1.53, 1.53, 
    1.53, 1.52, 1.51, 1.5, 1.49, 1.48, 1.47, 1.45, 1.44, 1.42, 1.41, 1.39, 
    1.38, 1.36, 1.35, 1.33, 1.32, 1.3, 1.29, 1.27, 1.26, 1.24, 1.23, 1.21, 
    1.2, 1.18, 1.16, 1.15, 1.13, 1.11, 1.09, 1.07, 1.05, 1.04, 1.02, 0.995, 
    0.974, 0.954, 0.933, 0.912, 0.891, 0.869, 0.848, 0.827, 0.807, 0.785, 
    0.764, 0.743, 0.722, 0.7, 0.679, 0.657, 0.635, 0.613, 0.591, 0.569, 
    0.548, 0.527, 0.507, 0.487, 0.468, 0.449, 0.432, 0.415, 0.399, 0.384, 
    0.369, 0.356, 0.343, 0.331, 0.319, 0.308, 0.298, 0.289, 0.28, 0.272, 
    0.265, 0.258, 0.252, 0.246, 0.241, 0.237, 0.233, 0.23, 0.227, 0.225, 
    0.223, 0.222, 0.221, 0.221, 0.22, 0.221, 0.221, 0.222, 0.222, 0.224, 
    0.225, 0.226, 0.228, 0.229, 0.231, 0.233, 0.235, 0.237, 0.239, 0.241, 
    0.244, 0.246, 0.248, 0.249, 0.251, 0.253, 0.255, 0.256, 0.257, 0.259, 
    0.259, 0.26, 0.26, 0.26, 0.259, 0.257, 0.255, 0.252, 0.248, 0.244, 0.239, 
    0.233, 0.227, 0.22, 0.214, 0.207, 0.2, 0.193, 0.187, 0.181, 0.175, 0.17, 
    0.165, 0.161, 0.158, 0.155, 0.153, 0.151, 0.149, 0.148, 0.147, 0.145, 
    0.144, 0.143, 0.142, 0.14, 0.139, 0.137, 0.136, 0.135, 0.133, 0.132, 
    0.13, 0.129, 0.128, 0.127, 0.126, 0.125, 0.124, 0.123, 0.122, 0.121, 
    0.12, 0.119, 0.119, 0.118, 0.117, 0.116, 0.116, 0.115, 0.115, 0.115, 
    0.114, 0.114, 0.114, 0.114, 0.113, 0.113, 0.113, 0.113, 0.113, 0.113, 
    0.113, 0.114, 0.115, 0.116, 0.117, 0.118, 0.12, 0.121, 0.122, 0.124, 
    0.125, 0.126, 0.126, 0.127, 0.127, 0.127, 0.126, 0.126, 0.125, 0.124, 
    0.123, 0.121, 0.12, 0.119, 0.117, 0.116, 0.114, 0.113, 0.112, 0.111, 
    0.111, 0.111, 0.112, 0.115, 0.119, 0.124, 0.131, 0.139, 0.148, 0.158, 
    0.169, 0.18, 0.191, 0.201, 0.211, 0.219, 0.225, 0.23, 0.232, 0.233, 
    0.231, 0.229, 0.226, 0.222, 0.218, 0.216, 0.214, 0.214, 0.215, 0.218, 
    0.221, 0.225, 0.23, 0.235, 0.239, 0.243, 0.245, 0.246, 0.246, 0.244, 
    0.241, 0.237, 0.233, 0.228, 0.223, 0.218, 0.213, 0.21, 0.207, 0.204, 
    0.203, 0.202, 0.202, 0.201, 0.202, 0.202, 0.203, 0.204, 0.204, 0.204, 
    0.205, 0.205, 0.205, 0.204, 0.203, 0.202, 0.201, 0.199, 0.197, 0.195, 
    0.193, 0.191, 0.188, 0.186, 0.184, 0.182, 0.18, 0.178, 0.177, 0.176, 
    0.175, 0.175, 0.174, 0.174, 0.174, 0.174, 0.174, 0.174, 0.174, 0.174, 
    0.173, 0.172, 0.172, 0.171, 0.17, 0.17, 0.169, 0.169, 0.168, 0.168, 
    0.168, 0.169, 0.169, 0.169, 0.169, 0.17, 0.171, 0.172, 0.173, 0.175, 
    0.176, 0.179, 0.181, 0.184, 0.188, 0.192, 0.196, 0.2, 0.203, 0.207, 0.21, 
    0.213, 0.215, 0.216, 0.216, 0.216, 0.216, 0.215, 0.213, 0.212, 0.21, 
    0.208, 0.207, 0.206, 0.205, 0.204, 0.203, 0.203, 0.203, 0.202, 0.202, 
    0.202, 0.201, 0.201, 0.201, 0.2, 0.199, 0.199, 0.198, 0.198, 0.198, 
    0.198, 0.197, 0.198, 0.198, 0.198, 0.199, 0.2, 0.201, 0.202, 0.203, 
    0.205, 0.206, 0.208, 0.21, 0.211, 0.213, 0.215, 0.217, 0.219, 0.221, 
    0.224, 0.226, 0.228, 0.23, 0.233, 0.235, 0.237, 0.24, 0.242, 0.245, 
    0.248, 0.25, 0.253, 0.256, 0.258, 0.261, 0.263, 0.265, 0.267, 0.269, 
    0.27, 0.271, 0.273, 0.274, 0.276, 0.278, 0.28, 0.282, 0.285, 0.288, 
    0.292, 0.296, 0.3, 0.304, 0.309, 0.313, 0.318, 0.324, 0.329, 0.335, 
    0.341, 0.347, 0.354, 0.361, 0.368, 0.376, 0.384, 0.392, 0.401, 0.41, 
    0.419, 0.429, 0.439, 0.449, 0.46, 0.471, 0.482, 0.493, 0.505, 0.516, 
    0.528, 0.54, 0.552, 0.565, 0.577, 0.59, 0.602, 0.615, 0.628, 0.64, 0.653, 
    0.666, 0.679, 0.692, 0.705, 0.719, 0.732, 0.746, 0.759, 0.773, 0.787, 
    0.8, 0.814, 0.828, 0.842, 0.856, 0.869, 0.883, 0.897, 0.911, 0.925, 0.94, 
    0.954, 0.969, 0.984, 1, 1.02, 1.03, 1.05, 1.06, 1.08, 1.1, 1.11, 1.12, 
    1.14, 1.15, 1.17, 1.18, 1.19, 1.2, 1.21, 1.21, 1.22, 1.22, 1.23, 1.23, 
    1.23, 1.23, 1.22, 1.22, 1.21, 1.21, 1.2, 1.19, 1.18, 1.18, 1.17, 1.15, 
    1.14, 1.13, 1.12, 1.11, 1.1, 1.09, 1.08, 1.07, 1.06, 1.06, 1.05, 1.05, 
    1.05, 1.05, 1.06, 1.06, 1.07, 1.08, 1.09, 1.1, 1.12, 1.13, 1.15, 1.17, 
    1.19, 1.21, 1.24, 1.26, 1.29, 1.32, 1.35, 1.38, 1.41, 1.44, 1.47, 1.5, 
    1.52, 1.55, 1.57, 1.59, 1.61, 1.62, 1.62, 1.63, 1.62, 1.61, 1.59, 1.57, 
    1.55, 1.52, 1.48, 1.45, 1.41, 1.37, 1.34, 1.3, 1.27, 1.23, 1.2, 1.18, 
    1.15, 1.12, 1.1, 1.08, 1.05, 1.03, 1.01, 0.984, 0.963, 0.942, 0.923, 
    0.906, 0.89, 0.877, 0.866, 0.857, 0.851, 0.846, 0.843, 0.842, 0.842, 
    0.842, 0.843, 0.844, 0.844, 0.844, 0.843, 0.84, 0.836, 0.83, 0.823, 
    0.814, 0.804, 0.791, 0.777, 0.762, 0.746, 0.729, 0.71, 0.691, 0.672, 
    0.652, 0.631, 0.61, 0.59, 0.57, 0.551, 0.535, 0.521, 0.51, 0.502, 0.499, 
    0.498, 0.501, 0.507, 0.515, 0.524, 0.533, 0.54, 0.546, 0.549, 0.548, 
    0.543, 0.534, 0.521, 0.506, 0.489, 0.472, 0.456, 0.441, 0.429, 0.421, 
    0.416, 0.414, 0.416, 0.422, 0.43, 0.44, 0.451, 0.463, 0.476, 0.488, 0.5, 
    0.51, 0.518, 0.524, 0.528, 0.529, 0.528, 0.525, 0.52, 0.514, 0.508, 
    0.501, 0.494, 0.488, 0.482, 0.477, 0.472, 0.468, 0.464, 0.459, 0.455, 
    0.449, 0.443, 0.436, 0.428, 0.419, 0.41, 0.4, 0.39, 0.379, 0.369, 0.359, 
    0.349, 0.34, 0.332, 0.324, 0.318, 0.312, 0.307, 0.303, 0.299, 0.296, 
    0.293, 0.29, 0.287, 0.284, 0.282, 0.279, 0.277, 0.274, 0.272, 0.27, 
    0.268, 0.265, 0.263, 0.261, 0.258, 0.256, 0.253, 0.25, 0.247, 0.244, 
    0.241, 0.239, 0.236, 0.233, 0.23, 0.228, 0.225, 0.222, 0.22, 0.218, 
    0.215, 0.213, 0.212, 0.21, 0.209, 0.208, 0.207, 0.206, 0.206, 0.206, 
    0.205, 0.205, 0.205, 0.205, 0.205, 0.205, 0.205, 0.206, 0.206, 0.206, 
    0.207, 0.208, 0.209, 0.21, 0.212, 0.214, 0.217, 0.221, 0.225, 0.23, 
    0.236, 0.242, 0.249, 0.256, 0.263, 0.27, 0.277, 0.283, 0.288, 0.292, 
    0.295, 0.297, 0.298, 0.298, 0.297, 0.295, 0.292, 0.288, 0.284, 0.279, 
    0.274, 0.268, 0.262, 0.256, 0.249, 0.242, 0.235, 0.228, 0.221, 0.214, 
    0.207, 0.201, 0.196, 0.191, 0.188, 0.185, 0.183, 0.18, 0.178, 0.177, 
    0.175, 0.173, 0.171, 0.169, 0.168, 0.167, 0.167, 0.167, 0.167, 0.166, 
    0.165, 0.164, 0.163, 0.162, 0.162, 0.162, 0.163, 0.164, 0.165, 0.165, 
    0.164, 0.164, 0.163, 0.162, 0.162, 0.162, 0.162, 0.163, 0.165, 0.167, 
    0.17, 0.172, 0.176, 0.18, 0.184, 0.188, 0.192, 0.196, 0.199, 0.202, 
    0.205, 0.208, 0.211, 0.214, 0.216, 0.218, 0.219, 0.219, 0.218, 0.216, 
    0.213, 0.209, 0.205, 0.201, 0.197, 0.193, 0.189, 0.186, 0.184, 0.181, 
    0.179, 0.177, 0.176, 0.175, 0.175, 0.176, 0.178, 0.18, 0.182, 0.185, 
    0.188, 0.191, 0.194, 0.196, 0.198, 0.198, 0.199, 0.2, 0.2, 0.201, 0.201, 
    0.202, 0.204, 0.206, 0.208, 0.21, 0.212, 0.215, 0.218, 0.22, 0.223, 
    0.227, 0.23, 0.234, 0.239, 0.244, 0.25, 0.255, 0.261, 0.266, 0.271, 
    0.274, 0.276, 0.278, 0.279, 0.28, 0.281, 0.281, 0.283, 0.284, 0.287, 
    0.29, 0.293, 0.296, 0.3, 0.305, 0.311, 0.318, 0.328, 0.34, 0.354, 0.368, 
    0.382, 0.395, 0.406, 0.415, 0.42, 0.423, 0.423, 0.421, 0.419, 0.416, 
    0.413, 0.409, 0.404, 0.398, 0.392, 0.386, 0.379, 0.37, 0.36, 0.349, 
    0.337, 0.325, 0.311, 0.297, 0.282, 0.267, 0.252, 0.235, 0.219, 0.201, 
    0.183, 0.166, 0.15, 0.136, 0.124, 0.113, 0.104, 0.097, 0.091, 0.086, 
    0.08, 0.075, 0.071, 0.068, 0.065, 0.064, 0.063, 0.062, 0.062, 0.062, 
    0.062, 0.061, 0.06, 0.059, 0.059, 0.059, 0.06, 0.061, 0.062, 0.063, 
    0.064, 0.066 ;

 bnd_kaolinite = 0.185, 0.19, 0.2, 0.21, 0.215, 0.22, 0.225, 0.233, 0.24, 0.26, 0.28, 
    0.3, 0.325, 0.36, 0.37, 0.4, 0.433, 0.466, 0.5, 0.533, 0.566, 0.6, 0.633, 
    0.666, 0.7, 0.817, 0.907, 1, 1.105, 1.2, 1.303, 1.4, 1.5, 1.6, 1.7, 1.8, 
    1.9, 2, 2.1, 2.2, 2.3, 2.4, 2.4999,
// NB: Relabel EgH79 value at 2.5 um as 2.4999 um to make room for 2.5 um Roush datum
// NB: Excise EgH79 value at 2.6 um in favor of Roush data
// end EgH79 Kaolinite. Begin Roush Kaolinite:
    2.5, 2.5006, 2.5013, 2.5019, 2.5025, 2.5031, 2.5038, 2.5044, 2.505, 
    2.5056, 2.5063, 2.5069, 2.5075, 2.5082, 2.5088, 2.5094, 2.51, 2.5107, 
    2.5113, 2.5119, 2.5126, 2.5132, 2.5138, 2.5145, 2.5151, 2.5157, 2.5164, 
    2.517, 2.5176, 2.5183, 2.5189, 2.5195, 2.5202, 2.5208, 2.5214, 2.5221, 
    2.5227, 2.5233, 2.524, 2.5246, 2.5253, 2.5259, 2.5265, 2.5272, 2.5278, 
    2.5284, 2.5291, 2.5297, 2.5304, 2.531, 2.5316, 2.5323, 2.5329, 2.5336, 
    2.5342, 2.5349, 2.5355, 2.5361, 2.5368, 2.5374, 2.5381, 2.5387, 2.5394, 
    2.54, 2.5407, 2.5413, 2.5419, 2.5426, 2.5432, 2.5439, 2.5445, 2.5452, 
    2.5458, 2.5465, 2.5471, 2.5478, 2.5484, 2.5491, 2.5497, 2.5504, 2.551, 
    2.5517, 2.5523, 2.553, 2.5536, 2.5543, 2.5549, 2.5556, 2.5562, 2.5569, 
    2.5575, 2.5582, 2.5589, 2.5595, 2.5602, 2.5608, 2.5615, 2.5621, 2.5628, 
    2.5634, 2.5641, 2.5648, 2.5654, 2.5661, 2.5667, 2.5674, 2.5681, 2.5687, 
    2.5694, 2.57, 2.5707, 2.5714, 2.572, 2.5727, 2.5733, 2.574, 2.5747, 
    2.5753, 2.576, 2.5767, 2.5773, 2.578, 2.5786, 2.5793, 2.58, 2.5806, 
    2.5813, 2.582, 2.5826, 2.5833, 2.584, 2.5846, 2.5853, 2.586, 2.5867, 
    2.5873, 2.588, 2.5887, 2.5893, 2.59, 2.5907, 2.5913, 2.592, 2.5927, 
    2.5934, 2.594, 2.5947, 2.5954, 2.5961, 2.5967, 2.5974, 2.5981, 2.5988, 
    2.5994, 2.6001, 2.6008, 2.6015, 2.6021, 2.6028, 2.6035, 2.6042, 2.6048, 
    2.6055, 2.6062, 2.6069, 2.6076, 2.6082, 2.6089, 2.6096, 2.6103, 2.611, 
    2.6116, 2.6123, 2.613, 2.6137, 2.6144, 2.6151, 2.6157, 2.6164, 2.6171, 
    2.6178, 2.6185, 2.6192, 2.6199, 2.6205, 2.6212, 2.6219, 2.6226, 2.6233, 
    2.624, 2.6247, 2.6254, 2.6261, 2.6267, 2.6274, 2.6281, 2.6288, 2.6295, 
    2.6302, 2.6309, 2.6316, 2.6323, 2.633, 2.6337, 2.6344, 2.635, 2.6357, 
    2.6364, 2.6371, 2.6378, 2.6385, 2.6392, 2.6399, 2.6406, 2.6413, 2.642, 
    2.6427, 2.6434, 2.6441, 2.6448, 2.6455, 2.6462, 2.6469, 2.6476, 2.6483, 
    2.649, 2.6497, 2.6504, 2.6511, 2.6518, 2.6525, 2.6532, 2.6539, 2.6546, 
    2.6553, 2.656, 2.6567, 2.6575, 2.6582, 2.6589, 2.6596, 2.6603, 2.661, 
    2.6617, 2.6624, 2.6631, 2.6638, 2.6645, 2.6652, 2.666, 2.6667, 2.6674, 
    2.6681, 2.6688, 2.6695, 2.6702, 2.6709, 2.6717, 2.6724, 2.6731, 2.6738, 
    2.6745, 2.6752, 2.6759, 2.6767, 2.6774, 2.6781, 2.6788, 2.6795, 2.6802, 
    2.681, 2.6817, 2.6824, 2.6831, 2.6838, 2.6846, 2.6853, 2.686, 2.6867, 
    2.6874, 2.6882, 2.6889, 2.6896, 2.6903, 2.6911, 2.6918, 2.6925, 2.6932, 
    2.694, 2.6947, 2.6954, 2.6961, 2.6969, 2.6976, 2.6983, 2.6991, 2.6998, 
    2.7005, 2.7012, 2.702, 2.7027, 2.7034, 2.7042, 2.7049, 2.7056, 2.7064, 
    2.7071, 2.7078, 2.7086, 2.7093, 2.71, 2.7108, 2.7115, 2.7122, 2.713, 
    2.7137, 2.7144, 2.7152, 2.7159, 2.7167, 2.7174, 2.7181, 2.7189, 2.7196, 
    2.7203, 2.7211, 2.7218, 2.7226, 2.7233, 2.7241, 2.7248, 2.7255, 2.7263, 
    2.727, 2.7278, 2.7285, 2.7293, 2.73, 2.7307, 2.7315, 2.7322, 2.733, 
    2.7337, 2.7345, 2.7352, 2.736, 2.7367, 2.7375, 2.7382, 2.739, 2.7397, 
    2.7405, 2.7412, 2.742, 2.7427, 2.7435, 2.7442, 2.745, 2.7457, 2.7465, 
    2.7473, 2.748, 2.7488, 2.7495, 2.7503, 2.751, 2.7518, 2.7525, 2.7533, 
    2.7541, 2.7548, 2.7556, 2.7563, 2.7571, 2.7579, 2.7586, 2.7594, 2.7601, 
    2.7609, 2.7617, 2.7624, 2.7632, 2.764, 2.7647, 2.7655, 2.7663, 2.767, 
    2.7678, 2.7685, 2.7693, 2.7701, 2.7709, 2.7716, 2.7724, 2.7732, 2.7739, 
    2.7747, 2.7755, 2.7762, 2.777, 2.7778, 2.7785, 2.7793, 2.7801, 2.7809, 
    2.7816, 2.7824, 2.7832, 2.784, 2.7847, 2.7855, 2.7863, 2.7871, 2.7878, 
    2.7886, 2.7894, 2.7902, 2.791, 2.7917, 2.7925, 2.7933, 2.7941, 2.7949, 
    2.7956, 2.7964, 2.7972, 2.798, 2.7988, 2.7996, 2.8003, 2.8011, 2.8019, 
    2.8027, 2.8035, 2.8043, 2.805, 2.8058, 2.8066, 2.8074, 2.8082, 2.809, 
    2.8098, 2.8106, 2.8114, 2.8121, 2.8129, 2.8137, 2.8145, 2.8153, 2.8161, 
    2.8169, 2.8177, 2.8185, 2.8193, 2.8201, 2.8209, 2.8217, 2.8225, 2.8233, 
    2.8241, 2.8249, 2.8257, 2.8265, 2.8273, 2.8281, 2.8289, 2.8297, 2.8305, 
    2.8313, 2.8321, 2.8329, 2.8337, 2.8345, 2.8353, 2.8361, 2.8369, 2.8377, 
    2.8385, 2.8393, 2.8401, 2.8409, 2.8417, 2.8425, 2.8433, 2.8441, 2.845, 
    2.8458, 2.8466, 2.8474, 2.8482, 2.849, 2.8498, 2.8506, 2.8514, 2.8523, 
    2.8531, 2.8539, 2.8547, 2.8555, 2.8563, 2.8571, 2.858, 2.8588, 2.8596, 
    2.8604, 2.8612, 2.862, 2.8629, 2.8637, 2.8645, 2.8653, 2.8662, 2.867, 
    2.8678, 2.8686, 2.8694, 2.8703, 2.8711, 2.8719, 2.8727, 2.8736, 2.8744, 
    2.8752, 2.876, 2.8769, 2.8777, 2.8785, 2.8794, 2.8802, 2.881, 2.8818, 
    2.8827, 2.8835, 2.8843, 2.8852, 2.886, 2.8868, 2.8877, 2.8885, 2.8893, 
    2.8902, 2.891, 2.8918, 2.8927, 2.8935, 2.8944, 2.8952, 2.896, 2.8969, 
    2.8977, 2.8986, 2.8994, 2.9002, 2.9011, 2.9019, 2.9028, 2.9036, 2.9044, 
    2.9053, 2.9061, 2.907, 2.9078, 2.9087, 2.9095, 2.9104, 2.9112, 2.9121, 
    2.9129, 2.9138, 2.9146, 2.9155, 2.9163, 2.9172, 2.918, 2.9189, 2.9197, 
    2.9206, 2.9214, 2.9223, 2.9231, 2.924, 2.9248, 2.9257, 2.9265, 2.9274, 
    2.9283, 2.9291, 2.93, 2.9308, 2.9317, 2.9326, 2.9334, 2.9343, 2.9351, 
    2.936, 2.9369, 2.9377, 2.9386, 2.9394, 2.9403, 2.9412, 2.942, 2.9429, 
    2.9438, 2.9446, 2.9455, 2.9464, 2.9472, 2.9481, 2.949, 2.9499, 2.9507, 
    2.9516, 2.9525, 2.9533, 2.9542, 2.9551, 2.956, 2.9568, 2.9577, 2.9586, 
    2.9595, 2.9603, 2.9612, 2.9621, 2.963, 2.9638, 2.9647, 2.9656, 2.9665, 
    2.9674, 2.9682, 2.9691, 2.97, 2.9709, 2.9718, 2.9727, 2.9735, 2.9744, 
    2.9753, 2.9762, 2.9771, 2.978, 2.9789, 2.9797, 2.9806, 2.9815, 2.9824, 
    2.9833, 2.9842, 2.9851, 2.986, 2.9869, 2.9878, 2.9886, 2.9895, 2.9904, 
    2.9913, 2.9922, 2.9931, 2.994, 2.9949, 2.9958, 2.9967, 2.9976, 2.9985, 
    2.9994, 3.0003, 3.0012, 3.0021, 3.003, 3.0039, 3.0048, 3.0057, 3.0066, 
    3.0075, 3.0084, 3.0093, 3.0102, 3.0111, 3.012, 3.013, 3.0139, 3.0148, 
    3.0157, 3.0166, 3.0175, 3.0184, 3.0193, 3.0202, 3.0211, 3.0221, 3.023, 
    3.0239, 3.0248, 3.0257, 3.0266, 3.0276, 3.0285, 3.0294, 3.0303, 3.0312, 
    3.0321, 3.0331, 3.034, 3.0349, 3.0358, 3.0367, 3.0377, 3.0386, 3.0395, 
    3.0404, 3.0414, 3.0423, 3.0432, 3.0441, 3.0451, 3.046, 3.0469, 3.0479, 
    3.0488, 3.0497, 3.0506, 3.0516, 3.0525, 3.0534, 3.0544, 3.0553, 3.0562, 
    3.0572, 3.0581, 3.059, 3.06, 3.0609, 3.0618, 3.0628, 3.0637, 3.0647, 
    3.0656, 3.0665, 3.0675, 3.0684, 3.0694, 3.0703, 3.0713, 3.0722, 3.0731, 
    3.0741, 3.075, 3.076, 3.0769, 3.0779, 3.0788, 3.0798, 3.0807, 3.0817, 
    3.0826, 3.0836, 3.0845, 3.0855, 3.0864, 3.0874, 3.0883, 3.0893, 3.0902, 
    3.0912, 3.0921, 3.0931, 3.0941, 3.095, 3.096, 3.0969, 3.0979, 3.0989, 
    3.0998, 3.1008, 3.1017, 3.1027, 3.1037, 3.1046, 3.1056, 3.1066, 3.1075, 
    3.1085, 3.1095, 3.1104, 3.1114, 3.1124, 3.1133, 3.1143, 3.1153, 3.1162, 
    3.1172, 3.1182, 3.1192, 3.1201, 3.1211, 3.1221, 3.123, 3.124, 3.125, 
    3.126, 3.127, 3.1279, 3.1289, 3.1299, 3.1309, 3.1319, 3.1328, 3.1338, 
    3.1348, 3.1358, 3.1368, 3.1377, 3.1387, 3.1397, 3.1407, 3.1417, 3.1427, 
    3.1437, 3.1447, 3.1456, 3.1466, 3.1476, 3.1486, 3.1496, 3.1506, 3.1516, 
    3.1526, 3.1536, 3.1546, 3.1556, 3.1566, 3.1576, 3.1586, 3.1596, 3.1606, 
    3.1616, 3.1626, 3.1636, 3.1646, 3.1656, 3.1666, 3.1676, 3.1686, 3.1696, 
    3.1706, 3.1716, 3.1726, 3.1736, 3.1746, 3.1756, 3.1766, 3.1776, 3.1786, 
    3.1797, 3.1807, 3.1817, 3.1827, 3.1837, 3.1847, 3.1857, 3.1867, 3.1878, 
    3.1888, 3.1898, 3.1908, 3.1918, 3.1928, 3.1939, 3.1949, 3.1959, 3.1969, 
    3.198, 3.199, 3.2, 3.201, 3.202, 3.2031, 3.2041, 3.2051, 3.2062, 3.2072, 
    3.2082, 3.2092, 3.2103, 3.2113, 3.2123, 3.2134, 3.2144, 3.2154, 3.2165, 
    3.2175, 3.2185, 3.2196, 3.2206, 3.2216, 3.2227, 3.2237, 3.2248, 3.2258, 
    3.2268, 3.2279, 3.2289, 3.23, 3.231, 3.2321, 3.2331, 3.2342, 3.2352, 
    3.2362, 3.2373, 3.2383, 3.2394, 3.2404, 3.2415, 3.2425, 3.2436, 3.2446, 
    3.2457, 3.2468, 3.2478, 3.2489, 3.2499, 3.251, 3.252, 3.2531, 3.2541, 
    3.2552, 3.2563, 3.2573, 3.2584, 3.2595, 3.2605, 3.2616, 3.2626, 3.2637, 
    3.2648, 3.2658, 3.2669, 3.268, 3.269, 3.2701, 3.2712, 3.2723, 3.2733, 
    3.2744, 3.2755, 3.2765, 3.2776, 3.2787, 3.2798, 3.2808, 3.2819, 3.283, 
    3.2841, 3.2852, 3.2862, 3.2873, 3.2884, 3.2895, 3.2906, 3.2916, 3.2927, 
    3.2938, 3.2949, 3.296, 3.2971, 3.2982, 3.2992, 3.3003, 3.3014, 3.3025, 
    3.3036, 3.3047, 3.3058, 3.3069, 3.308, 3.3091, 3.3102, 3.3113, 3.3124, 
    3.3135, 3.3146, 3.3156, 3.3167, 3.3179, 3.319, 3.3201, 3.3212, 3.3223, 
    3.3234, 3.3245, 3.3256, 3.3267, 3.3278, 3.3289, 3.33, 3.3311, 3.3322, 
    3.3333, 3.3344, 3.3356, 3.3367, 3.3378, 3.3389, 3.34, 3.3411, 3.3422, 
    3.3434, 3.3445, 3.3456, 3.3467, 3.3478, 3.349, 3.3501, 3.3512, 3.3523, 
    3.3535, 3.3546, 3.3557, 3.3568, 3.358, 3.3591, 3.3602, 3.3613, 3.3625, 
    3.3636, 3.3647, 3.3659, 3.367, 3.3681, 3.3693, 3.3704, 3.3715, 3.3727, 
    3.3738, 3.375, 3.3761, 3.3772, 3.3784, 3.3795, 3.3807, 3.3818, 3.3829, 
    3.3841, 3.3852, 3.3864, 3.3875, 3.3887, 3.3898, 3.391, 3.3921, 3.3933, 
    3.3944, 3.3956, 3.3967, 3.3979, 3.399, 3.4002, 3.4014, 3.4025, 3.4037, 
    3.4048, 3.406, 3.4072, 3.4083, 3.4095, 3.4106, 3.4118, 3.413, 3.4141, 
    3.4153, 3.4165, 3.4176, 3.4188, 3.42, 3.4211, 3.4223, 3.4235, 3.4247, 
    3.4258, 3.427, 3.4282, 3.4294, 3.4305, 3.4317, 3.4329, 3.4341, 3.4352, 
    3.4364, 3.4376, 3.4388, 3.44, 3.4412, 3.4423, 3.4435, 3.4447, 3.4459, 
    3.4471, 3.4483, 3.4495, 3.4507, 3.4518, 3.453, 3.4542, 3.4554, 3.4566, 
    3.4578, 3.459, 3.4602, 3.4614, 3.4626, 3.4638, 3.465, 3.4662, 3.4674, 
    3.4686, 3.4698, 3.471, 3.4722, 3.4734, 3.4746, 3.4758, 3.4771, 3.4783, 
    3.4795, 3.4807, 3.4819, 3.4831, 3.4843, 3.4855, 3.4868, 3.488, 3.4892, 
    3.4904, 3.4916, 3.4928, 3.4941, 3.4953, 3.4965, 3.4977, 3.499, 3.5002, 
    3.5014, 3.5026, 3.5039, 3.5051, 3.5063, 3.5075, 3.5088, 3.51, 3.5112, 
    3.5125, 3.5137, 3.5149, 3.5162, 3.5174, 3.5186, 3.5199, 3.5211, 3.5224, 
    3.5236, 3.5249, 3.5261, 3.5273, 3.5286, 3.5298, 3.5311, 3.5323, 3.5336, 
    3.5348, 3.5361, 3.5373, 3.5386, 3.5398, 3.5411, 3.5423, 3.5436, 3.5448, 
    3.5461, 3.5474, 3.5486, 3.5499, 3.5511, 3.5524, 3.5537, 3.5549, 3.5562, 
    3.5575, 3.5587, 3.56, 3.5613, 3.5625, 3.5638, 3.5651, 3.5663, 3.5676, 
    3.5689, 3.5702, 3.5714, 3.5727, 3.574, 3.5753, 3.5765, 3.5778, 3.5791, 
    3.5804, 3.5817, 3.5829, 3.5842, 3.5855, 3.5868, 3.5881, 3.5894, 3.5907, 
    3.592, 3.5932, 3.5945, 3.5958, 3.5971, 3.5984, 3.5997, 3.601, 3.6023, 
    3.6036, 3.6049, 3.6062, 3.6075, 3.6088, 3.6101, 3.6114, 3.6127, 3.614, 
    3.6153, 3.6166, 3.6179, 3.6193, 3.6206, 3.6219, 3.6232, 3.6245, 3.6258, 
    3.6271, 3.6284, 3.6298, 3.6311, 3.6324, 3.6337, 3.635, 3.6364, 3.6377, 
    3.639, 3.6403, 3.6417, 3.643, 3.6443, 3.6456, 3.647, 3.6483, 3.6496, 
    3.651, 3.6523, 3.6536, 3.655, 3.6563, 3.6576, 3.659, 3.6603, 3.6617, 
    3.663, 3.6643, 3.6657, 3.667, 3.6684, 3.6697, 3.6711, 3.6724, 3.6738, 
    3.6751, 3.6765, 3.6778, 3.6792, 3.6805, 3.6819, 3.6832, 3.6846, 3.686, 
    3.6873, 3.6887, 3.69, 3.6914, 3.6928, 3.6941, 3.6955, 3.6969, 3.6982, 
    3.6996, 3.701, 3.7023, 3.7037, 3.7051, 3.7064, 3.7078, 3.7092, 3.7106, 
    3.712, 3.7133, 3.7147, 3.7161, 3.7175, 3.7189, 3.7202, 3.7216, 3.723, 
    3.7244, 3.7258, 3.7272, 3.7286, 3.73, 3.7313, 3.7327, 3.7341, 3.7355, 
    3.7369, 3.7383, 3.7397, 3.7411, 3.7425, 3.7439, 3.7453, 3.7467, 3.7481, 
    3.7495, 3.7509, 3.7523, 3.7538, 3.7552, 3.7566, 3.758, 3.7594, 3.7608, 
    3.7622, 3.7636, 3.7651, 3.7665, 3.7679, 3.7693, 3.7707, 3.7722, 3.7736, 
    3.775, 3.7764, 3.7779, 3.7793, 3.7807, 3.7821, 3.7836, 3.785, 3.7864, 
    3.7879, 3.7893, 3.7908, 3.7922, 3.7936, 3.7951, 3.7965, 3.7979, 3.7994, 
    3.8008, 3.8023, 3.8037, 3.8052, 3.8066, 3.8081, 3.8095, 3.811, 3.8124, 
    3.8139, 3.8153, 3.8168, 3.8183, 3.8197, 3.8212, 3.8226, 3.8241, 3.8256, 
    3.827, 3.8285, 3.83, 3.8314, 3.8329, 3.8344, 3.8358, 3.8373, 3.8388, 
    3.8402, 3.8417, 3.8432, 3.8447, 3.8462, 3.8476, 3.8491, 3.8506, 3.8521, 
    3.8536, 3.8551, 3.8565, 3.858, 3.8595, 3.861, 3.8625, 3.864, 3.8655, 
    3.867, 3.8685, 3.87, 3.8715, 3.873, 3.8745, 3.876, 3.8775, 3.879, 3.8805, 
    3.882, 3.8835, 3.885, 3.8865, 3.888, 3.8895, 3.8911, 3.8926, 3.8941, 
    3.8956, 3.8971, 3.8986, 3.9002, 3.9017, 3.9032, 3.9047, 3.9063, 3.9078, 
    3.9093, 3.9108, 3.9124, 3.9139, 3.9154, 3.917, 3.9185, 3.92, 3.9216, 
    3.9231, 3.9246, 3.9262, 3.9277, 3.9293, 3.9308, 3.9324, 3.9339, 3.9355, 
    3.937, 3.9386, 3.9401, 3.9417, 3.9432, 3.9448, 3.9463, 3.9479, 3.9494, 
    3.951, 3.9526, 3.9541, 3.9557, 3.9573, 3.9588, 3.9604, 3.962, 3.9635, 
    3.9651, 3.9667, 3.9683, 3.9698, 3.9714, 3.973, 3.9746, 3.9761, 3.9777, 
    3.9793, 3.9809, 3.9825, 3.9841, 3.9857, 3.9872, 3.9888, 3.9904, 3.992, 
    3.9936, 3.9952, 3.9968, 3.9984, 4, 4.0016, 4.0032, 4.0048, 4.0064, 4.008, 
    4.0096, 4.0112, 4.0128, 4.0145, 4.0161, 4.0177, 4.0193, 4.0209, 4.0225, 
    4.0241, 4.0258, 4.0274, 4.029, 4.0306, 4.0323, 4.0339, 4.0355, 4.0371, 
    4.0388, 4.0404, 4.042, 4.0437, 4.0453, 4.0469, 4.0486, 4.0502, 4.0519, 
    4.0535, 4.0552, 4.0568, 4.0584, 4.0601, 4.0617, 4.0634, 4.065, 4.0667, 
    4.0683, 4.07, 4.0717, 4.0733, 4.075, 4.0766, 4.0783, 4.08, 4.0816, 
    4.0833, 4.085, 4.0866, 4.0883, 4.09, 4.0917, 4.0933, 4.095, 4.0967, 
    4.0984, 4.1, 4.1017, 4.1034, 4.1051, 4.1068, 4.1085, 4.1102, 4.1118, 
    4.1135, 4.1152, 4.1169, 4.1186, 4.1203, 4.122, 4.1237, 4.1254, 4.1271, 
    4.1288, 4.1305, 4.1322, 4.1339, 4.1356, 4.1374, 4.1391, 4.1408, 4.1425, 
    4.1442, 4.1459, 4.1477, 4.1494, 4.1511, 4.1528, 4.1545, 4.1563, 4.158, 
    4.1597, 4.1615, 4.1632, 4.1649, 4.1667, 4.1684, 4.1701, 4.1719, 4.1736, 
    4.1754, 4.1771, 4.1789, 4.1806, 4.1824, 4.1841, 4.1859, 4.1876, 4.1894, 
    4.1911, 4.1929, 4.1946, 4.1964, 4.1982, 4.1999, 4.2017, 4.2034, 4.2052, 
    4.207, 4.2088, 4.2105, 4.2123, 4.2141, 4.2159, 4.2176, 4.2194, 4.2212, 
    4.223, 4.2248, 4.2265, 4.2283, 4.2301, 4.2319, 4.2337, 4.2355, 4.2373, 
    4.2391, 4.2409, 4.2427, 4.2445, 4.2463, 4.2481, 4.2499, 4.2517, 4.2535, 
    4.2553, 4.2571, 4.2589, 4.2608, 4.2626, 4.2644, 4.2662, 4.268, 4.2699, 
    4.2717, 4.2735, 4.2753, 4.2772, 4.279, 4.2808, 4.2827, 4.2845, 4.2863, 
    4.2882, 4.29, 4.2918, 4.2937, 4.2955, 4.2974, 4.2992, 4.3011, 4.3029, 
    4.3048, 4.3066, 4.3085, 4.3103, 4.3122, 4.3141, 4.3159, 4.3178, 4.3197, 
    4.3215, 4.3234, 4.3253, 4.3271, 4.329, 4.3309, 4.3328, 4.3346, 4.3365, 
    4.3384, 4.3403, 4.3422, 4.344, 4.3459, 4.3478, 4.3497, 4.3516, 4.3535, 
    4.3554, 4.3573, 4.3592, 4.3611, 4.363, 4.3649, 4.3668, 4.3687, 4.3706, 
    4.3725, 4.3745, 4.3764, 4.3783, 4.3802, 4.3821, 4.384, 4.386, 4.3879, 
    4.3898, 4.3917, 4.3937, 4.3956, 4.3975, 4.3995, 4.4014, 4.4033, 4.4053, 
    4.4072, 4.4092, 4.4111, 4.4131, 4.415, 4.417, 4.4189, 4.4209, 4.4228, 
    4.4248, 4.4267, 4.4287, 4.4307, 4.4326, 4.4346, 4.4366, 4.4385, 4.4405, 
    4.4425, 4.4444, 4.4464, 4.4484, 4.4504, 4.4524, 4.4543, 4.4563, 4.4583, 
    4.4603, 4.4623, 4.4643, 4.4663, 4.4683, 4.4703, 4.4723, 4.4743, 4.4763, 
    4.4783, 4.4803, 4.4823, 4.4843, 4.4863, 4.4883, 4.4903, 4.4924, 4.4944, 
    4.4964, 4.4984, 4.5005, 4.5025, 4.5045, 4.5065, 4.5086, 4.5106, 4.5126, 
    4.5147, 4.5167, 4.5188, 4.5208, 4.5228, 4.5249, 4.5269, 4.529, 4.531, 
    4.5331, 4.5351, 4.5372, 4.5393, 4.5413, 4.5434, 4.5455, 4.5475, 4.5496, 
    4.5517, 4.5537, 4.5558, 4.5579, 4.56, 4.562, 4.5641, 4.5662, 4.5683, 
    4.5704, 4.5725, 4.5746, 4.5767, 4.5788, 4.5809, 4.583, 4.5851, 4.5872, 
    4.5893, 4.5914, 4.5935, 4.5956, 4.5977, 4.5998, 4.6019, 4.6041, 4.6062, 
    4.6083, 4.6104, 4.6125, 4.6147, 4.6168, 4.6189, 4.6211, 4.6232, 4.6253, 
    4.6275, 4.6296, 4.6318, 4.6339, 4.6361, 4.6382, 4.6404, 4.6425, 4.6447, 
    4.6468, 4.649, 4.6512, 4.6533, 4.6555, 4.6577, 4.6598, 4.662, 4.6642, 
    4.6664, 4.6685, 4.6707, 4.6729, 4.6751, 4.6773, 4.6795, 4.6816, 4.6838, 
    4.686, 4.6882, 4.6904, 4.6926, 4.6948, 4.697, 4.6992, 4.7015, 4.7037, 
    4.7059, 4.7081, 4.7103, 4.7125, 4.7148, 4.717, 4.7192, 4.7214, 4.7237, 
    4.7259, 4.7281, 4.7304, 4.7326, 4.7348, 4.7371, 4.7393, 4.7416, 4.7438, 
    4.7461, 4.7483, 4.7506, 4.7529, 4.7551, 4.7574, 4.7596, 4.7619, 4.7642, 
    4.7664, 4.7687, 4.771, 4.7733, 4.7755, 4.7778, 4.7801, 4.7824, 4.7847, 
    4.787, 4.7893, 4.7916, 4.7939, 4.7962, 4.7985, 4.8008, 4.8031, 4.8054, 
    4.8077, 4.81, 4.8123, 4.8146, 4.817, 4.8193, 4.8216, 4.8239, 4.8263, 
    4.8286, 4.8309, 4.8333, 4.8356, 4.8379, 4.8403, 4.8426, 4.845, 4.8473, 
    4.8497, 4.852, 4.8544, 4.8567, 4.8591, 4.8614, 4.8638, 4.8662, 4.8685, 
    4.8709, 4.8733, 4.8757, 4.878, 4.8804, 4.8828, 4.8852, 4.8876, 4.89, 
    4.8924, 4.8948, 4.8972, 4.8996, 4.902, 4.9044, 4.9068, 4.9092, 4.9116, 
    4.914, 4.9164, 4.9188, 4.9213, 4.9237, 4.9261, 4.9285, 4.931, 4.9334, 
    4.9358, 4.9383, 4.9407, 4.9432, 4.9456, 4.948, 4.9505, 4.9529, 4.9554, 
    4.9579, 4.9603, 4.9628, 4.9652, 4.9677, 4.9702, 4.9727, 4.9751, 4.9776, 
    4.9801, 4.9826, 4.985, 4.9875, 4.99, 4.9925, 4.995, 4.9975, 5, 5.0025, 
    5.005, 5.0075, 5.01, 5.0125, 5.015, 5.0176, 5.0201, 5.0226, 5.0251, 
    5.0277, 5.0302, 5.0327, 5.0352, 5.0378, 5.0403, 5.0429, 5.0454, 5.048, 
    5.0505, 5.0531, 5.0556, 5.0582, 5.0607, 5.0633, 5.0659, 5.0684, 5.071, 
    5.0736, 5.0761, 5.0787, 5.0813, 5.0839, 5.0865, 5.0891, 5.0916, 5.0942, 
    5.0968, 5.0994, 5.102, 5.1046, 5.1073, 5.1099, 5.1125, 5.1151, 5.1177, 
    5.1203, 5.123, 5.1256, 5.1282, 5.1308, 5.1335, 5.1361, 5.1387, 5.1414, 
    5.144, 5.1467, 5.1493, 5.152, 5.1546, 5.1573, 5.16, 5.1626, 5.1653, 
    5.168, 5.1706, 5.1733, 5.176, 5.1787, 5.1813, 5.184, 5.1867, 5.1894, 
    5.1921, 5.1948, 5.1975, 5.2002, 5.2029, 5.2056, 5.2083, 5.211, 5.2138, 
    5.2165, 5.2192, 5.2219, 5.2247, 5.2274, 5.2301, 5.2329, 5.2356, 5.2383, 
    5.2411, 5.2438, 5.2466, 5.2493, 5.2521, 5.2549, 5.2576, 5.2604, 5.2632, 
    5.2659, 5.2687, 5.2715, 5.2743, 5.277, 5.2798, 5.2826, 5.2854, 5.2882, 
    5.291, 5.2938, 5.2966, 5.2994, 5.3022, 5.305, 5.3079, 5.3107, 5.3135, 
    5.3163, 5.3191, 5.322, 5.3248, 5.3277, 5.3305, 5.3333, 5.3362, 5.339, 
    5.3419, 5.3447, 5.3476, 5.3505, 5.3533, 5.3562, 5.3591, 5.3619, 5.3648, 
    5.3677, 5.3706, 5.3735, 5.3763, 5.3792, 5.3821, 5.385, 5.3879, 5.3908, 
    5.3937, 5.3967, 5.3996, 5.4025, 5.4054, 5.4083, 5.4113, 5.4142, 5.4171, 
    5.4201, 5.423, 5.4259, 5.4289, 5.4318, 5.4348, 5.4377, 5.4407, 5.4437, 
    5.4466, 5.4496, 5.4526, 5.4555, 5.4585, 5.4615, 5.4645, 5.4675, 5.4705, 
    5.4735, 5.4765, 5.4795, 5.4825, 5.4855, 5.4885, 5.4915, 5.4945, 5.4975, 
    5.5006, 5.5036, 5.5066, 5.5096, 5.5127, 5.5157, 5.5188, 5.5218, 5.5249, 
    5.5279, 5.531, 5.534, 5.5371, 5.5402, 5.5432, 5.5463, 5.5494, 5.5525, 
    5.5556, 5.5586, 5.5617, 5.5648, 5.5679, 5.571, 5.5741, 5.5772, 5.5804, 
    5.5835, 5.5866, 5.5897, 5.5928, 5.596, 5.5991, 5.6022, 5.6054, 5.6085, 
    5.6117, 5.6148, 5.618, 5.6211, 5.6243, 5.6275, 5.6306, 5.6338, 5.637, 
    5.6402, 5.6433, 5.6465, 5.6497, 5.6529, 5.6561, 5.6593, 5.6625, 5.6657, 
    5.6689, 5.6721, 5.6754, 5.6786, 5.6818, 5.685, 5.6883, 5.6915, 5.6948, 
    5.698, 5.7013, 5.7045, 5.7078, 5.711, 5.7143, 5.7176, 5.7208, 5.7241, 
    5.7274, 5.7307, 5.7339, 5.7372, 5.7405, 5.7438, 5.7471, 5.7504, 5.7537, 
    5.7571, 5.7604, 5.7637, 5.767, 5.7703, 5.7737, 5.777, 5.7803, 5.7837, 
    5.787, 5.7904, 5.7937, 5.7971, 5.8005, 5.8038, 5.8072, 5.8106, 5.814, 
    5.8173, 5.8207, 5.8241, 5.8275, 5.8309, 5.8343, 5.8377, 5.8411, 5.8445, 
    5.848, 5.8514, 5.8548, 5.8582, 5.8617, 5.8651, 5.8685, 5.872, 5.8754, 
    5.8789, 5.8824, 5.8858, 5.8893, 5.8928, 5.8962, 5.8997, 5.9032, 5.9067, 
    5.9102, 5.9137, 5.9172, 5.9207, 5.9242, 5.9277, 5.9312, 5.9347, 5.9382, 
    5.9418, 5.9453, 5.9488, 5.9524, 5.9559, 5.9595, 5.963, 5.9666, 5.9701, 
    5.9737, 5.9773, 5.9809, 5.9844, 5.988, 5.9916, 5.9952, 5.9988, 6.0024, 
    6.006, 6.0096, 6.0132, 6.0168, 6.0205, 6.0241, 6.0277, 6.0314, 6.035, 
    6.0386, 6.0423, 6.0459, 6.0496, 6.0533, 6.0569, 6.0606, 6.0643, 6.068, 
    6.0716, 6.0753, 6.079, 6.0827, 6.0864, 6.0901, 6.0938, 6.0976, 6.1013, 
    6.105, 6.1087, 6.1125, 6.1162, 6.12, 6.1237, 6.1275, 6.1312, 6.135, 
    6.1387, 6.1425, 6.1463, 6.1501, 6.1538, 6.1576, 6.1614, 6.1652, 6.169, 
    6.1728, 6.1767, 6.1805, 6.1843, 6.1881, 6.192, 6.1958, 6.1996, 6.2035, 
    6.2073, 6.2112, 6.215, 6.2189, 6.2228, 6.2267, 6.2305, 6.2344, 6.2383, 
    6.2422, 6.2461, 6.25, 6.2539, 6.2578, 6.2617, 6.2657, 6.2696, 6.2735, 
    6.2775, 6.2814, 6.2854, 6.2893, 6.2933, 6.2972, 6.3012, 6.3052, 6.3091, 
    6.3131, 6.3171, 6.3211, 6.3251, 6.3291, 6.3331, 6.3371, 6.3412, 6.3452, 
    6.3492, 6.3532, 6.3573, 6.3613, 6.3654, 6.3694, 6.3735, 6.3776, 6.3816, 
    6.3857, 6.3898, 6.3939, 6.398, 6.402, 6.4061, 6.4103, 6.4144, 6.4185, 
    6.4226, 6.4267, 6.4309, 6.435, 6.4392, 6.4433, 6.4475, 6.4516, 6.4558, 
    6.4599, 6.4641, 6.4683, 6.4725, 6.4767, 6.4809, 6.4851, 6.4893, 6.4935, 
    6.4977, 6.502, 6.5062, 6.5104, 6.5147, 6.5189, 6.5232, 6.5274, 6.5317, 
    6.5359, 6.5402, 6.5445, 6.5488, 6.5531, 6.5574, 6.5617, 6.566, 6.5703, 
    6.5746, 6.5789, 6.5833, 6.5876, 6.592, 6.5963, 6.6007, 6.605, 6.6094, 
    6.6138, 6.6181, 6.6225, 6.6269, 6.6313, 6.6357, 6.6401, 6.6445, 6.6489, 
    6.6534, 6.6578, 6.6622, 6.6667, 6.6711, 6.6756, 6.68, 6.6845, 6.689, 
    6.6934, 6.6979, 6.7024, 6.7069, 6.7114, 6.7159, 6.7204, 6.7249, 6.7295, 
    6.734, 6.7385, 6.7431, 6.7476, 6.7522, 6.7568, 6.7613, 6.7659, 6.7705, 
    6.7751, 6.7797, 6.7843, 6.7889, 6.7935, 6.7981, 6.8027, 6.8074, 6.812, 
    6.8166, 6.8213, 6.8259, 6.8306, 6.8353, 6.8399, 6.8446, 6.8493, 6.854, 
    6.8587, 6.8634, 6.8681, 6.8729, 6.8776, 6.8823, 6.8871, 6.8918, 6.8966, 
    6.9013, 6.9061, 6.9109, 6.9156, 6.9204, 6.9252, 6.93, 6.9348, 6.9396, 
    6.9444, 6.9493, 6.9541, 6.9589, 6.9638, 6.9686, 6.9735, 6.9784, 6.9832, 
    6.9881, 6.993, 6.9979, 7.0028, 7.0077, 7.0126, 7.0175, 7.0225, 7.0274, 
    7.0323, 7.0373, 7.0423, 7.0472, 7.0522, 7.0572, 7.0621, 7.0671, 7.0721, 
    7.0771, 7.0822, 7.0872, 7.0922, 7.0972, 7.1023, 7.1073, 7.1124, 7.1174, 
    7.1225, 7.1276, 7.1327, 7.1378, 7.1429, 7.148, 7.1531, 7.1582, 7.1633, 
    7.1685, 7.1736, 7.1788, 7.1839, 7.1891, 7.1942, 7.1994, 7.2046, 7.2098, 
    7.215, 7.2202, 7.2254, 7.2307, 7.2359, 7.2411, 7.2464, 7.2516, 7.2569, 
    7.2622, 7.2674, 7.2727, 7.278, 7.2833, 7.2886, 7.2939, 7.2993, 7.3046, 
    7.3099, 7.3153, 7.3206, 7.326, 7.3314, 7.3368, 7.3421, 7.3475, 7.3529, 
    7.3584, 7.3638, 7.3692, 7.3746, 7.3801, 7.3855, 7.391, 7.3964, 7.4019, 
    7.4074, 7.4129, 7.4184, 7.4239, 7.4294, 7.4349, 7.4405, 7.446, 7.4516, 
    7.4571, 7.4627, 7.4683, 7.4738, 7.4794, 7.485, 7.4906, 7.4963, 7.5019, 
    7.5075, 7.5131, 7.5188, 7.5245, 7.5301, 7.5358, 7.5415, 7.5472, 7.5529, 
    7.5586, 7.5643, 7.57, 7.5758, 7.5815, 7.5873, 7.593, 7.5988, 7.6046, 
    7.6104, 7.6161, 7.622, 7.6278, 7.6336, 7.6394, 7.6453, 7.6511, 7.657, 
    7.6628, 7.6687, 7.6746, 7.6805, 7.6864, 7.6923, 7.6982, 7.7042, 7.7101, 
    7.716, 7.722, 7.728, 7.734, 7.7399, 7.7459, 7.7519, 7.758, 7.764, 7.77, 
    7.776, 7.7821, 7.7882, 7.7942, 7.8003, 7.8064, 7.8125, 7.8186, 7.8247, 
    7.8309, 7.837, 7.8431, 7.8493, 7.8555, 7.8616, 7.8678, 7.874, 7.8802, 
    7.8864, 7.8927, 7.8989, 7.9051, 7.9114, 7.9177, 7.9239, 7.9302, 7.9365, 
    7.9428, 7.9491, 7.9554, 7.9618, 7.9681, 7.9745, 7.9808, 7.9872, 7.9936, 
    8, 8.0064, 8.0128, 8.0192, 8.0257, 8.0321, 8.0386, 8.0451, 8.0515, 8.058, 
    8.0645, 8.071, 8.0775, 8.0841, 8.0906, 8.0972, 8.1037, 8.1103, 8.1169, 
    8.1235, 8.1301, 8.1367, 8.1433, 8.15, 8.1566, 8.1633, 8.1699, 8.1766, 
    8.1833, 8.19, 8.1967, 8.2034, 8.2102, 8.2169, 8.2237, 8.2305, 8.2372, 
    8.244, 8.2508, 8.2576, 8.2645, 8.2713, 8.2781, 8.285, 8.2919, 8.2988, 
    8.3056, 8.3126, 8.3195, 8.3264, 8.3333, 8.3403, 8.3472, 8.3542, 8.3612, 
    8.3682, 8.3752, 8.3822, 8.3893, 8.3963, 8.4034, 8.4104, 8.4175, 8.4246, 
    8.4317, 8.4388, 8.4459, 8.4531, 8.4602, 8.4674, 8.4746, 8.4818, 8.489, 
    8.4962, 8.5034, 8.5106, 8.5179, 8.5251, 8.5324, 8.5397, 8.547, 8.5543, 
    8.5616, 8.569, 8.5763, 8.5837, 8.5911, 8.5985, 8.6059, 8.6133, 8.6207, 
    8.6281, 8.6356, 8.643, 8.6505, 8.658, 8.6655, 8.673, 8.6806, 8.6881, 
    8.6957, 8.7032, 8.7108, 8.7184, 8.726, 8.7336, 8.7413, 8.7489, 8.7566, 
    8.7642, 8.7719, 8.7796, 8.7873, 8.7951, 8.8028, 8.8106, 8.8183, 8.8261, 
    8.8339, 8.8417, 8.8496, 8.8574, 8.8652, 8.8731, 8.881, 8.8889, 8.8968, 
    8.9047, 8.9127, 8.9206, 8.9286, 8.9366, 8.9445, 8.9526, 8.9606, 8.9686, 
    8.9767, 8.9847, 8.9928, 9.0009, 9.009, 9.0171, 9.0253, 9.0334, 9.0416, 
    9.0498, 9.058, 9.0662, 9.0744, 9.0827, 9.0909, 9.0992, 9.1075, 9.1158, 
    9.1241, 9.1324, 9.1408, 9.1491, 9.1575, 9.1659, 9.1743, 9.1827, 9.1912, 
    9.1996, 9.2081, 9.2166, 9.2251, 9.2336, 9.2421, 9.2507, 9.2593, 9.2678, 
    9.2764, 9.2851, 9.2937, 9.3023, 9.311, 9.3197, 9.3284, 9.3371, 9.3458, 
    9.3545, 9.3633, 9.3721, 9.3809, 9.3897, 9.3985, 9.4073, 9.4162, 9.4251, 
    9.434, 9.4429, 9.4518, 9.4607, 9.4697, 9.4787, 9.4877, 9.4967, 9.5057, 
    9.5147, 9.5238, 9.5329, 9.542, 9.5511, 9.5602, 9.5694, 9.5785, 9.5877, 
    9.5969, 9.6061, 9.6154, 9.6246, 9.6339, 9.6432, 9.6525, 9.6618, 9.6712, 
    9.6805, 9.6899, 9.6993, 9.7087, 9.7182, 9.7276, 9.7371, 9.7466, 9.7561, 
    9.7656, 9.7752, 9.7847, 9.7943, 9.8039, 9.8135, 9.8232, 9.8328, 9.8425, 
    9.8522, 9.8619, 9.8717, 9.8814, 9.8912, 9.901, 9.9108, 9.9206, 9.9305, 
    9.9404, 9.9502, 9.9602, 9.9701, 9.98, 9.99, 10, 10.01, 10.02, 10.03, 
    10.04, 10.05, 10.06, 10.071, 10.081, 10.091, 10.101, 10.111, 10.122, 
    10.132, 10.142, 10.152, 10.163, 10.173, 10.183, 10.194, 10.204, 10.215, 
    10.225, 10.235, 10.246, 10.256, 10.267, 10.278, 10.288, 10.299, 10.309, 
    10.32, 10.331, 10.341, 10.352, 10.363, 10.373, 10.384, 10.395, 10.406, 
    10.417, 10.427, 10.438, 10.449, 10.46, 10.471, 10.482, 10.493, 10.504, 
    10.515, 10.526, 10.537, 10.549, 10.56, 10.571, 10.582, 10.593, 10.604, 
    10.616, 10.627, 10.638, 10.65, 10.661, 10.672, 10.684, 10.695, 10.707, 
    10.718, 10.73, 10.741, 10.753, 10.764, 10.776, 10.788, 10.799, 10.811, 
    10.823, 10.834, 10.846, 10.858, 10.87, 10.881, 10.893, 10.905, 10.917, 
    10.929, 10.941, 10.953, 10.965, 10.977, 10.989, 11.001, 11.013, 11.025, 
    11.038, 11.05, 11.062, 11.074, 11.087, 11.099, 11.111, 11.123, 11.136, 
    11.148, 11.161, 11.173, 11.186, 11.198, 11.211, 11.223, 11.236, 11.249, 
    11.261, 11.274, 11.287, 11.299, 11.312, 11.325, 11.338, 11.351, 11.364, 
    11.377, 11.389, 11.403, 11.415, 11.429, 11.442, 11.455, 11.468, 11.481, 
    11.494, 11.507, 11.521, 11.534, 11.547, 11.561, 11.574, 11.587, 11.601, 
    11.614, 11.628, 11.641, 11.655, 11.669, 11.682, 11.696, 11.71, 11.723, 
    11.737, 11.751, 11.765, 11.779, 11.792, 11.806, 11.82, 11.834, 11.848, 
    11.862, 11.877, 11.891, 11.905, 11.919, 11.933, 11.947, 11.962, 11.976, 
    11.99, 12.005, 12.019, 12.034, 12.048, 12.063, 12.077, 12.092, 12.106, 
    12.121, 12.136, 12.151, 12.165, 12.18, 12.195, 12.21, 12.225, 12.24, 
    12.255, 12.27, 12.285, 12.3, 12.315, 12.33, 12.346, 12.361, 12.376, 
    12.392, 12.407, 12.422, 12.438, 12.453, 12.469, 12.484, 12.5, 12.516, 
    12.531, 12.547, 12.563, 12.579, 12.594, 12.61, 12.626, 12.642, 12.658, 
    12.674, 12.69, 12.707, 12.723, 12.739, 12.755, 12.771, 12.788, 12.804, 
    12.821, 12.837, 12.854, 12.87, 12.887, 12.903, 12.92, 12.937, 12.953, 
    12.97, 12.987, 13.004, 13.021, 13.038, 13.055, 13.072, 13.089, 13.106, 
    13.123, 13.141, 13.158, 13.175, 13.193, 13.21, 13.227, 13.245, 13.263, 
    13.28, 13.298, 13.316, 13.333, 13.351, 13.369, 13.387, 13.405, 13.423, 
    13.441, 13.459, 13.477, 13.495, 13.514, 13.532, 13.55, 13.568, 13.587, 
    13.605, 13.624, 13.643, 13.661, 13.68, 13.699, 13.717, 13.736, 13.755, 
    13.774, 13.793, 13.812, 13.831, 13.85, 13.87, 13.889, 13.908, 13.928, 
    13.947, 13.967, 13.986, 14.006, 14.025, 14.045, 14.065, 14.085, 14.104, 
    14.124, 14.144, 14.164, 14.184, 14.205, 14.225, 14.245, 14.265, 14.286, 
    14.306, 14.327, 14.347, 14.368, 14.389, 14.409, 14.43, 14.451, 14.472, 
    14.493, 14.514, 14.535, 14.556, 14.577, 14.599, 14.62, 14.641, 14.663, 
    14.684, 14.706, 14.727, 14.749, 14.771, 14.793, 14.815, 14.837, 14.859, 
    14.881, 14.903, 14.925, 14.948, 14.97, 14.993, 15.015, 15.038, 15.06, 
    15.083, 15.106, 15.129, 15.151, 15.175, 15.198, 15.221, 15.244, 15.267, 
    15.29, 15.314, 15.337, 15.361, 15.385, 15.408, 15.432, 15.456, 15.48, 
    15.504, 15.528, 15.552, 15.576, 15.601, 15.625, 15.649, 15.674, 15.699, 
    15.723, 15.748, 15.773, 15.798, 15.823, 15.848, 15.873, 15.898, 15.924, 
    15.949, 15.974, 16, 16.026, 16.051, 16.077, 16.103, 16.129, 16.155, 
    16.181, 16.208, 16.234, 16.26, 16.287, 16.313, 16.34, 16.367, 16.393, 
    16.42, 16.447, 16.475, 16.502, 16.529, 16.556, 16.584, 16.611, 16.639, 
    16.667, 16.694, 16.722, 16.75, 16.778, 16.807, 16.835, 16.863, 16.892, 
    16.92, 16.949, 16.978, 17.007, 17.036, 17.065, 17.094, 17.123, 17.153, 
    17.182, 17.212, 17.241, 17.271, 17.301, 17.331, 17.361, 17.391, 17.422, 
    17.452, 17.483, 17.513, 17.544, 17.575, 17.606, 17.637, 17.668, 17.699, 
    17.73, 17.762, 17.794, 17.825, 17.857, 17.889, 17.921, 17.953, 17.986, 
    18.018, 18.051, 18.083, 18.116, 18.149, 18.182, 18.215, 18.248, 18.281, 
    18.315, 18.349, 18.382, 18.416, 18.45, 18.484, 18.518, 18.553, 18.587, 
    18.622, 18.657, 18.692, 18.727, 18.762, 18.797, 18.832, 18.868, 18.904, 
    18.939, 18.975, 19.011, 19.048, 19.084, 19.121, 19.157, 19.194, 19.231, 
    19.268, 19.305, 19.342, 19.38, 19.417, 19.455, 19.493, 19.531, 19.569, 
    19.608, 19.646, 19.685, 19.724, 19.763, 19.802, 19.841, 19.881, 19.92, 
    19.96, 20, 20.04, 20.08, 20.121, 20.161, 20.202, 20.243, 20.284, 20.325, 
    20.367, 20.408, 20.45, 20.492, 20.534, 20.576, 20.619, 20.661, 20.704, 
    20.747, 20.79, 20.833, 20.877, 20.92, 20.964, 21.008, 21.053, 21.097, 
    21.142, 21.186, 21.231, 21.277, 21.322, 21.368, 21.413, 21.459, 21.505, 
    21.552, 21.598, 21.645, 21.692, 21.739, 21.787, 21.834, 21.882, 21.93, 
    21.978, 22.026, 22.075, 22.124, 22.173, 22.222, 22.272, 22.321, 22.371, 
    22.421, 22.472, 22.522, 22.573, 22.624, 22.676, 22.727, 22.779, 22.831, 
    22.883, 22.936, 22.989, 23.042, 23.095, 23.148, 23.202, 23.256, 23.31, 
    23.365, 23.419, 23.474, 23.529, 23.585, 23.641, 23.697, 23.753, 23.809, 
    23.866, 23.923, 23.981, 24.038, 24.096, 24.155, 24.213, 24.272, 24.331, 
    24.39, 24.45, 24.51, 24.57, 24.631, 24.691, 24.753, 24.814, 24.876, 
    24.938, 25, 25.063, 25.126, 25.189, 25.253, 25.316, 25.381, 25.445, 
    25.51, 25.575, 25.641, 25.707, 25.773, 25.84, 25.907, 25.974, 26.042, 
    26.11, 26.178, 26.247, 26.316, 26.385, 26.455, 26.525, 26.596, 26.667, 
    26.738, 26.81, 26.882, 26.954, 27.027, 27.1, 27.174, 27.248, 27.322, 
    27.397, 27.472, 27.548, 27.624, 27.701, 27.778, 27.855, 27.933, 28.011, 
    28.09, 28.169, 28.249, 28.329, 28.409, 28.49, 28.571, 28.653, 28.736, 
    28.818, 28.902, 28.986, 29.07, 29.154, 29.24, 29.326, 29.412, 29.499, 
    29.586, 29.674, 29.762, 29.851, 29.94, 30.03, 30.121, 30.212, 30.303, 
    30.395, 30.488, 30.581, 30.675, 30.769, 30.864, 30.96, 31.056, 31.153, 
    31.25, 31.348, 31.447, 31.546, 31.646, 31.746, 31.847, 31.949, 32.051, 
    32.154, 32.258, 32.362, 32.467, 32.573, 32.68, 32.787, 32.895, 33.003, 
    33.113, 33.223, 33.333, 33.445, 33.557, 33.67, 33.784, 33.898, 34.014, 
    34.13, 34.247, 34.364, 34.483, 34.602, 34.722, 34.843, 34.965, 35.088, 
    35.211, 35.336, 35.461, 35.587, 35.714, 35.842, 35.971, 36.101, 36.232, 
    36.364, 36.496, 36.63, 36.765, 36.9, 37.037, 37.175, 37.313, 37.453, 
    37.594, 37.736, 37.879, 38.023, 38.168, 38.314, 38.461, 38.61, 38.76, 
    38.91, 39.062, 39.216, 39.37, 39.526, 39.682, 39.841, 40, 40.161, 40.323, 
    40.486, 40.65, 40.816, 40.984, 41.152, 41.322, 41.494, 41.667, 41.841, 
    42.017, 42.194, 42.373, 42.553, 42.735, 42.918, 43.103, 43.29, 43.478, 
    43.668, 43.86, 44.053, 44.248, 44.444, 44.643, 44.843, 45.045, 45.249, 
    45.454, 45.662, 45.872, 46.083, 46.296, 46.512, 46.729, 46.948, 47.17, 
    47.393, 47.619, 47.847, 48.077, 48.309, 48.544, 48.78, 49.02, 49.261, 
    49.505, 49.751, 50, 50.251, 50.505, 50.761, 51.02, 51.282, 51.546, 
    51.813, 52.083, 52.356, 52.632, 52.91, 53.192, 53.476, 53.763, 54.054, 
    54.348, 54.645, 54.945, 55.249, 55.556, 55.866, 56.18, 56.497, 56.818, 
    57.143, 57.471, 57.804, 58.139, 58.479, 58.824, 59.172, 59.524, 59.88, 
    60.241, 60.606, 60.976, 61.35, 61.728, 62.112, 62.5, 62.893, 63.291, 
    63.694, 64.103, 64.516, 64.935, 65.359, 65.789, 66.225, 66.667, 67.114, 
    67.568, 68.027, 68.493, 68.965, 69.444, 69.93, 70.423, 70.922, 71.429, 
    71.942, 72.464, 72.993, 73.529, 74.074, 74.627, 75.188, 75.758, 76.336, 
    76.923, 77.519, 78.125, 78.74, 79.365, 80, 80.645, 81.301, 81.967, 
    82.645, 83.333, 84.034, 84.746, 85.47, 86.207, 86.956, 87.719, 88.496, 
    89.286, 90.09, 90.909, 91.743, 92.593, 93.458, 94.34, 95.238, 96.154, 
    97.087, 98.039, 99.01, 100, 101.01, 102.04, 103.09, 104.17, 105.26, 
    106.38, 107.53, 108.7, 109.89, 111.11, 112.36, 113.64, 114.94, 116.28, 
    117.65, 119.05, 120.48, 121.95, 123.46, 125, 126.58, 128.21, 129.87, 
    131.58, 133.33, 135.14, 136.99, 138.89, 140.85, 142.86, 144.93, 147.06, 
    149.25, 151.52, 153.85, 156.25, 158.73, 161.29, 163.93, 166.67, 169.49, 
    172.41, 175.44, 178.57, 181.82, 185.19, 188.68, 192.31, 196.08, 200 ;

 idx_rfr_kaolinite_rl = 1.491, 1.494, 1.496, 1.498, 1.501, 1.503, 1.506, 
    1.508, 1.511, 1.513, 1.506, 1.514, 1.512, 1.509, 1.5, 1.49, 1.491, 1.492, 
    1.493, 1.493, 1.493, 1.493, 1.494, 1.496, 1.497, 1.499, 1.501, 1.502, 
    1.502, 1.502, 1.502, 1.502, 1.502, 1.502, 1.502, 1.502, 1.502, 1.502, 
    1.502, 1.502, 1.502, 1.502, 1.502,
// NB: Relabel EgH79 value at 2.5 um as 2.4999 um to make room for 2.5 um Roush datum
// NB: Excise EgH79 value at 2.6 um in favor of Roush data
// end EgH79 Kaolinite. Begin Roush Kaolinite:
    1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 
    1.362, 1.362, 1.361, 1.361, 1.361, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 
    1.36, 1.361, 1.361, 1.362, 1.362, 1.363, 1.363, 1.363, 1.363, 1.362, 
    1.362, 1.361, 1.361, 1.36, 1.36, 1.36, 1.359, 1.359, 1.36, 1.36, 1.36, 
    1.361, 1.361, 1.362, 1.362, 1.362, 1.362, 1.362, 1.363, 1.363, 1.363, 
    1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.362, 1.362, 
    1.361, 1.361, 1.36, 1.36, 1.36, 1.36, 1.361, 1.361, 1.361, 1.362, 1.362, 
    1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.362, 
    1.361, 1.361, 1.36, 1.36, 1.359, 1.359, 1.359, 1.359, 1.359, 1.36, 1.36, 
    1.361, 1.361, 1.361, 1.362, 1.362, 1.361, 1.361, 1.361, 1.36, 1.36, 1.36, 
    1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.359, 1.359, 1.358, 
    1.358, 1.358, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.358, 
    1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 
    1.357, 1.357, 1.357, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.359, 
    1.359, 1.359, 1.359, 1.358, 1.358, 1.358, 1.358, 1.358, 1.359, 1.359, 
    1.359, 1.36, 1.36, 1.361, 1.361, 1.361, 1.361, 1.361, 1.36, 1.359, 1.358, 
    1.358, 1.357, 1.356, 1.356, 1.355, 1.355, 1.355, 1.356, 1.356, 1.356, 
    1.357, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.357, 1.357, 1.357, 
    1.357, 1.356, 1.356, 1.356, 1.357, 1.357, 1.358, 1.358, 1.359, 1.359, 
    1.36, 1.36, 1.36, 1.36, 1.359, 1.359, 1.359, 1.358, 1.358, 1.358, 1.358, 
    1.357, 1.357, 1.357, 1.356, 1.356, 1.355, 1.355, 1.355, 1.354, 1.354, 
    1.353, 1.353, 1.353, 1.353, 1.353, 1.353, 1.353, 1.352, 1.352, 1.352, 
    1.352, 1.351, 1.351, 1.351, 1.35, 1.35, 1.35, 1.35, 1.35, 1.35, 1.35, 
    1.35, 1.35, 1.35, 1.35, 1.349, 1.349, 1.349, 1.349, 1.349, 1.348, 1.348, 
    1.348, 1.348, 1.348, 1.349, 1.349, 1.349, 1.349, 1.348, 1.348, 1.348, 
    1.347, 1.346, 1.344, 1.343, 1.342, 1.341, 1.339, 1.338, 1.337, 1.336, 
    1.336, 1.335, 1.335, 1.336, 1.336, 1.336, 1.336, 1.336, 1.336, 1.335, 
    1.334, 1.333, 1.332, 1.33, 1.328, 1.326, 1.324, 1.322, 1.32, 1.318, 
    1.316, 1.314, 1.313, 1.311, 1.31, 1.308, 1.307, 1.306, 1.305, 1.304, 
    1.304, 1.304, 1.305, 1.306, 1.307, 1.309, 1.311, 1.314, 1.317, 1.32, 
    1.324, 1.327, 1.33, 1.333, 1.335, 1.337, 1.339, 1.341, 1.342, 1.343, 
    1.345, 1.345, 1.346, 1.346, 1.347, 1.347, 1.347, 1.347, 1.347, 1.347, 
    1.346, 1.346, 1.346, 1.346, 1.345, 1.346, 1.346, 1.346, 1.347, 1.347, 
    1.348, 1.348, 1.349, 1.35, 1.35, 1.351, 1.351, 1.352, 1.352, 1.353, 
    1.353, 1.354, 1.354, 1.355, 1.355, 1.355, 1.355, 1.355, 1.356, 1.356, 
    1.355, 1.355, 1.354, 1.353, 1.352, 1.351, 1.349, 1.347, 1.345, 1.343, 
    1.34, 1.338, 1.335, 1.334, 1.334, 1.334, 1.337, 1.341, 1.347, 1.355, 
    1.364, 1.374, 1.385, 1.396, 1.406, 1.415, 1.423, 1.429, 1.432, 1.434, 
    1.433, 1.431, 1.427, 1.424, 1.419, 1.415, 1.411, 1.407, 1.404, 1.402, 
    1.4, 1.398, 1.397, 1.397, 1.396, 1.396, 1.396, 1.396, 1.396, 1.395, 
    1.395, 1.395, 1.395, 1.394, 1.393, 1.392, 1.392, 1.391, 1.39, 1.389, 
    1.388, 1.387, 1.386, 1.386, 1.385, 1.385, 1.385, 1.384, 1.384, 1.384, 
    1.384, 1.383, 1.383, 1.383, 1.382, 1.382, 1.381, 1.381, 1.38, 1.38, 1.38, 
    1.379, 1.379, 1.379, 1.379, 1.379, 1.38, 1.38, 1.38, 1.38, 1.38, 1.381, 
    1.381, 1.381, 1.381, 1.381, 1.381, 1.381, 1.38, 1.38, 1.38, 1.379, 1.379, 
    1.379, 1.379, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.378, 1.378, 1.377, 
    1.377, 1.377, 1.376, 1.376, 1.376, 1.375, 1.375, 1.375, 1.375, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.375, 1.375, 1.375, 1.375, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.373, 1.373, 1.373, 1.373, 1.373, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 
    1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 
    1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.378, 1.378, 1.378, 1.378, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 1.376, 
    1.376, 1.376, 1.376, 1.376, 1.376, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.372, 
    1.372, 1.372, 1.372, 1.373, 1.373, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.364, 1.364, 
    1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 
    1.364, 1.364, 1.364, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 
    1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.362, 1.362, 
    1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 
    1.362, 1.362, 1.362, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 
    1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 
    1.361, 1.361, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 
    1.36, 1.36, 1.36, 1.36, 1.36, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 
    1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.358, 
    1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 
    1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 
    1.358, 1.358, 1.358, 1.358, 1.358, 1.357, 1.357, 1.357, 1.357, 1.357, 
    1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 
    1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 
    1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 
    1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 
    1.356, 1.356, 1.356, 1.356, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 
    1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 
    1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 
    1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 
    1.355, 1.355, 1.355, 1.355, 1.354, 1.354, 1.354, 1.354, 1.354, 1.354, 
    1.354, 1.354, 1.354, 1.354, 1.354, 1.354, 1.354, 1.354, 1.354, 1.354, 
    1.354, 1.354, 1.354, 1.354, 1.354, 1.354, 1.354, 1.354, 1.354, 1.353, 
    1.353, 1.353, 1.353, 1.353, 1.353, 1.353, 1.353, 1.353, 1.353, 1.353, 
    1.353, 1.353, 1.353, 1.353, 1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 
    1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 
    1.352, 1.352, 1.352, 1.352, 1.351, 1.351, 1.351, 1.351, 1.351, 1.351, 
    1.351, 1.351, 1.351, 1.351, 1.351, 1.351, 1.351, 1.351, 1.351, 1.35, 
    1.35, 1.35, 1.35, 1.35, 1.35, 1.35, 1.35, 1.35, 1.35, 1.35, 1.35, 1.35, 
    1.35, 1.35, 1.349, 1.349, 1.349, 1.349, 1.349, 1.349, 1.349, 1.349, 
    1.349, 1.349, 1.349, 1.349, 1.349, 1.349, 1.349, 1.348, 1.348, 1.348, 
    1.348, 1.348, 1.348, 1.348, 1.348, 1.348, 1.348, 1.347, 1.347, 1.347, 
    1.347, 1.347, 1.347, 1.347, 1.347, 1.347, 1.347, 1.347, 1.347, 1.347, 
    1.347, 1.347, 1.346, 1.346, 1.346, 1.346, 1.346, 1.346, 1.346, 1.346, 
    1.346, 1.346, 1.346, 1.346, 1.345, 1.345, 1.346, 1.345, 1.345, 1.345, 
    1.345, 1.345, 1.345, 1.345, 1.345, 1.345, 1.345, 1.344, 1.344, 1.344, 
    1.344, 1.344, 1.344, 1.344, 1.344, 1.344, 1.343, 1.343, 1.343, 1.343, 
    1.343, 1.343, 1.342, 1.342, 1.342, 1.342, 1.342, 1.342, 1.342, 1.342, 
    1.342, 1.342, 1.341, 1.341, 1.341, 1.341, 1.341, 1.341, 1.341, 1.34, 
    1.34, 1.34, 1.34, 1.34, 1.34, 1.34, 1.34, 1.34, 1.339, 1.339, 1.34, 
    1.339, 1.339, 1.339, 1.339, 1.339, 1.339, 1.338, 1.338, 1.338, 1.338, 
    1.338, 1.338, 1.338, 1.338, 1.338, 1.337, 1.337, 1.337, 1.337, 1.337, 
    1.337, 1.336, 1.336, 1.336, 1.336, 1.336, 1.336, 1.336, 1.336, 1.336, 
    1.335, 1.335, 1.335, 1.335, 1.335, 1.335, 1.335, 1.334, 1.334, 1.334, 
    1.334, 1.334, 1.334, 1.333, 1.333, 1.333, 1.333, 1.333, 1.333, 1.333, 
    1.332, 1.332, 1.332, 1.332, 1.332, 1.332, 1.332, 1.331, 1.331, 1.331, 
    1.331, 1.331, 1.331, 1.33, 1.33, 1.33, 1.33, 1.33, 1.33, 1.33, 1.329, 
    1.329, 1.329, 1.329, 1.329, 1.329, 1.328, 1.328, 1.328, 1.328, 1.328, 
    1.327, 1.327, 1.327, 1.327, 1.327, 1.326, 1.326, 1.326, 1.326, 1.326, 
    1.325, 1.325, 1.325, 1.325, 1.325, 1.324, 1.324, 1.324, 1.324, 1.324, 
    1.323, 1.323, 1.323, 1.323, 1.323, 1.322, 1.322, 1.322, 1.322, 1.322, 
    1.322, 1.322, 1.321, 1.321, 1.321, 1.321, 1.321, 1.32, 1.321, 1.32, 1.32, 
    1.32, 1.32, 1.319, 1.32, 1.319, 1.319, 1.319, 1.319, 1.319, 1.318, 1.318, 
    1.318, 1.318, 1.318, 1.317, 1.317, 1.317, 1.317, 1.317, 1.317, 1.317, 
    1.316, 1.316, 1.316, 1.316, 1.316, 1.315, 1.315, 1.315, 1.315, 1.315, 
    1.314, 1.314, 1.314, 1.314, 1.314, 1.313, 1.313, 1.313, 1.312, 1.313, 
    1.312, 1.312, 1.312, 1.312, 1.312, 1.311, 1.311, 1.311, 1.311, 1.311, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.309, 1.309, 1.309, 1.309, 1.308, 1.308, 
    1.308, 1.308, 1.307, 1.307, 1.307, 1.307, 1.306, 1.306, 1.306, 1.305, 
    1.305, 1.305, 1.305, 1.304, 1.304, 1.304, 1.304, 1.303, 1.303, 1.303, 
    1.303, 1.303, 1.302, 1.302, 1.302, 1.302, 1.301, 1.301, 1.301, 1.301, 
    1.3, 1.3, 1.3, 1.3, 1.299, 1.299, 1.299, 1.299, 1.298, 1.298, 1.298, 
    1.298, 1.297, 1.297, 1.297, 1.297, 1.296, 1.296, 1.296, 1.296, 1.295, 
    1.295, 1.295, 1.294, 1.294, 1.294, 1.294, 1.293, 1.293, 1.293, 1.293, 
    1.292, 1.292, 1.292, 1.292, 1.291, 1.291, 1.291, 1.291, 1.29, 1.29, 1.29, 
    1.289, 1.289, 1.289, 1.288, 1.288, 1.287, 1.287, 1.287, 1.286, 1.286, 
    1.286, 1.285, 1.285, 1.285, 1.284, 1.284, 1.284, 1.283, 1.283, 1.283, 
    1.282, 1.282, 1.282, 1.281, 1.281, 1.281, 1.28, 1.28, 1.28, 1.279, 1.279, 
    1.279, 1.278, 1.278, 1.277, 1.276, 1.276, 1.276, 1.275, 1.275, 1.275, 
    1.274, 1.274, 1.274, 1.273, 1.273, 1.272, 1.272, 1.272, 1.271, 1.27, 
    1.27, 1.27, 1.269, 1.269, 1.269, 1.268, 1.268, 1.268, 1.267, 1.266, 
    1.266, 1.266, 1.265, 1.265, 1.264, 1.264, 1.264, 1.263, 1.263, 1.262, 
    1.262, 1.262, 1.261, 1.261, 1.26, 1.26, 1.26, 1.259, 1.259, 1.258, 1.258, 
    1.257, 1.257, 1.256, 1.256, 1.256, 1.255, 1.254, 1.254, 1.254, 1.254, 
    1.253, 1.253, 1.252, 1.252, 1.251, 1.25, 1.25, 1.249, 1.249, 1.249, 
    1.248, 1.247, 1.247, 1.246, 1.246, 1.246, 1.245, 1.245, 1.244, 1.244, 
    1.243, 1.243, 1.242, 1.242, 1.241, 1.24, 1.24, 1.239, 1.239, 1.238, 
    1.237, 1.237, 1.236, 1.235, 1.235, 1.235, 1.234, 1.234, 1.233, 1.233, 
    1.232, 1.231, 1.231, 1.23, 1.229, 1.229, 1.228, 1.228, 1.227, 1.226, 
    1.226, 1.225, 1.224, 1.224, 1.224, 1.223, 1.222, 1.222, 1.221, 1.221, 
    1.22, 1.219, 1.219, 1.218, 1.217, 1.216, 1.215, 1.215, 1.214, 1.213, 
    1.213, 1.212, 1.212, 1.211, 1.21, 1.21, 1.209, 1.208, 1.207, 1.206, 
    1.206, 1.205, 1.204, 1.203, 1.202, 1.202, 1.201, 1.2, 1.2, 1.199, 1.198, 
    1.197, 1.196, 1.195, 1.194, 1.193, 1.192, 1.191, 1.19, 1.188, 1.187, 
    1.186, 1.185, 1.184, 1.182, 1.181, 1.18, 1.179, 1.178, 1.177, 1.177, 
    1.176, 1.175, 1.174, 1.173, 1.172, 1.171, 1.171, 1.17, 1.169, 1.168, 
    1.167, 1.167, 1.166, 1.165, 1.165, 1.164, 1.163, 1.162, 1.161, 1.161, 
    1.16, 1.159, 1.159, 1.158, 1.157, 1.156, 1.155, 1.154, 1.153, 1.152, 
    1.151, 1.149, 1.148, 1.147, 1.146, 1.145, 1.144, 1.143, 1.141, 1.14, 
    1.139, 1.138, 1.137, 1.135, 1.135, 1.133, 1.132, 1.13, 1.129, 1.127, 
    1.126, 1.124, 1.123, 1.121, 1.12, 1.118, 1.117, 1.115, 1.113, 1.112, 
    1.11, 1.109, 1.107, 1.106, 1.105, 1.103, 1.102, 1.1, 1.099, 1.097, 1.095, 
    1.094, 1.092, 1.091, 1.089, 1.087, 1.086, 1.084, 1.082, 1.081, 1.079, 
    1.077, 1.076, 1.074, 1.072, 1.071, 1.069, 1.067, 1.065, 1.063, 1.061, 
    1.059, 1.057, 1.055, 1.053, 1.051, 1.049, 1.046, 1.044, 1.041, 1.038, 
    1.035, 1.033, 1.03, 1.028, 1.025, 1.022, 1.02, 1.017, 1.015, 1.012, 1.01, 
    1.008, 1.005, 1.003, 1.001, 0.998, 0.995, 0.993, 0.99, 0.988, 0.985, 
    0.982, 0.98, 0.977, 0.974, 0.971, 0.967, 0.964, 0.961, 0.957, 0.953, 
    0.95, 0.946, 0.942, 0.938, 0.935, 0.931, 0.927, 0.923, 0.919, 0.914, 
    0.91, 0.906, 0.901, 0.897, 0.892, 0.887, 0.883, 0.878, 0.873, 0.868, 
    0.863, 0.857, 0.852, 0.847, 0.841, 0.836, 0.83, 0.825, 0.819, 0.812, 
    0.806, 0.8, 0.792, 0.785, 0.777, 0.769, 0.759, 0.75, 0.74, 0.729, 0.718, 
    0.707, 0.695, 0.683, 0.67, 0.658, 0.645, 0.633, 0.621, 0.608, 0.597, 
    0.585, 0.574, 0.564, 0.554, 0.545, 0.536, 0.529, 0.522, 0.516, 0.512, 
    0.508, 0.506, 0.505, 0.506, 0.509, 0.513, 0.518, 0.526, 0.535, 0.546, 
    0.56, 0.574, 0.591, 0.609, 0.629, 0.649, 0.67, 0.69, 0.71, 0.729, 0.746, 
    0.761, 0.772, 0.781, 0.786, 0.787, 0.784, 0.778, 0.769, 0.757, 0.743, 
    0.727, 0.709, 0.689, 0.669, 0.649, 0.628, 0.608, 0.587, 0.567, 0.548, 
    0.529, 0.511, 0.494, 0.478, 0.463, 0.449, 0.436, 0.424, 0.413, 0.404, 
    0.395, 0.388, 0.382, 0.377, 0.374, 0.371, 0.37, 0.37, 0.371, 0.372, 
    0.375, 0.379, 0.384, 0.389, 0.395, 0.403, 0.411, 0.419, 0.429, 0.439, 
    0.45, 0.462, 0.475, 0.489, 0.503, 0.519, 0.535, 0.553, 0.572, 0.592, 
    0.614, 0.637, 0.662, 0.689, 0.719, 0.751, 0.787, 0.826, 0.869, 0.917, 
    0.97, 1.028, 1.093, 1.164, 1.241, 1.324, 1.413, 1.506, 1.602, 1.699, 
    1.796, 1.888, 1.976, 2.055, 2.125, 2.184, 2.234, 2.273, 2.302, 2.324, 
    2.338, 2.346, 2.35, 2.351, 2.35, 2.347, 2.344, 2.341, 2.34, 2.339, 2.34, 
    2.343, 2.348, 2.356, 2.367, 2.382, 2.4, 2.421, 2.446, 2.475, 2.506, 2.54, 
    2.576, 2.613, 2.649, 2.684, 2.715, 2.741, 2.76, 2.77, 2.771, 2.762, 
    2.744, 2.716, 2.68, 2.638, 2.591, 2.541, 2.49, 2.438, 2.388, 2.339, 
    2.293, 2.249, 2.209, 2.171, 2.136, 2.104, 2.073, 2.045, 2.018, 1.993, 
    1.968, 1.945, 1.921, 1.899, 1.877, 1.855, 1.833, 1.812, 1.791, 1.77, 
    1.751, 1.732, 1.713, 1.696, 1.679, 1.663, 1.649, 1.636, 1.624, 1.613, 
    1.603, 1.595, 1.587, 1.581, 1.575, 1.57, 1.566, 1.562, 1.559, 1.556, 
    1.554, 1.552, 1.551, 1.55, 1.549, 1.549, 1.55, 1.552, 1.555, 1.558, 
    1.563, 1.569, 1.577, 1.586, 1.596, 1.609, 1.623, 1.638, 1.656, 1.675, 
    1.695, 1.717, 1.74, 1.764, 1.789, 1.815, 1.842, 1.869, 1.897, 1.926, 
    1.955, 1.983, 2.012, 2.04, 2.067, 2.093, 2.116, 2.138, 2.156, 2.172, 
    2.184, 2.192, 2.196, 2.196, 2.192, 2.185, 2.174, 2.161, 2.145, 2.128, 
    2.109, 2.089, 2.069, 2.049, 2.03, 2.011, 1.994, 1.977, 1.961, 1.946, 
    1.933, 1.921, 1.909, 1.898, 1.888, 1.878, 1.869, 1.86, 1.851, 1.843, 
    1.835, 1.827, 1.819, 1.811, 1.803, 1.796, 1.789, 1.782, 1.775, 1.768, 
    1.761, 1.755, 1.748, 1.742, 1.735, 1.729, 1.723, 1.717, 1.711, 1.705, 
    1.699, 1.694, 1.688, 1.683, 1.677, 1.672, 1.667, 1.662, 1.656, 1.651, 
    1.646, 1.641, 1.636, 1.631, 1.626, 1.621, 1.616, 1.611, 1.606, 1.601, 
    1.596, 1.591, 1.586, 1.581, 1.576, 1.571, 1.565, 1.56, 1.555, 1.549, 
    1.544, 1.538, 1.532, 1.526, 1.52, 1.514, 1.508, 1.502, 1.497, 1.491, 
    1.486, 1.481, 1.476, 1.472, 1.468, 1.465, 1.461, 1.459, 1.457, 1.455, 
    1.453, 1.452, 1.452, 1.452, 1.452, 1.453, 1.454, 1.455, 1.456, 1.458, 
    1.46, 1.462, 1.464, 1.466, 1.468, 1.47, 1.472, 1.474, 1.475, 1.476, 
    1.477, 1.477, 1.477, 1.476, 1.475, 1.473, 1.471, 1.468, 1.465, 1.461, 
    1.457, 1.452, 1.448, 1.443, 1.438, 1.433, 1.428, 1.423, 1.419, 1.414, 
    1.41, 1.406, 1.402, 1.398, 1.395, 1.392, 1.389, 1.387, 1.385, 1.383, 
    1.381, 1.379, 1.378, 1.377, 1.375, 1.374, 1.373, 1.372, 1.371, 1.37, 
    1.369, 1.368, 1.366, 1.365, 1.363, 1.361, 1.359, 1.357, 1.354, 1.351, 
    1.348, 1.344, 1.339, 1.335, 1.33, 1.324, 1.319, 1.312, 1.306, 1.3, 1.293, 
    1.285, 1.278, 1.271, 1.263, 1.256, 1.248, 1.241, 1.234, 1.227, 1.22, 
    1.214, 1.207, 1.201, 1.195, 1.19, 1.184, 1.179, 1.174, 1.17, 1.165, 
    1.161, 1.157, 1.154, 1.15, 1.147, 1.145, 1.142, 1.14, 1.138, 1.137, 
    1.135, 1.134, 1.132, 1.131, 1.13, 1.128, 1.127, 1.126, 1.125, 1.123, 
    1.122, 1.12, 1.118, 1.116, 1.114, 1.111, 1.108, 1.105, 1.102, 1.098, 
    1.094, 1.09, 1.086, 1.082, 1.077, 1.072, 1.067, 1.063, 1.057, 1.052, 
    1.047, 1.042, 1.038, 1.033, 1.028, 1.023, 1.019, 1.014, 1.01, 1.006, 
    1.002, 0.997, 0.993, 0.988, 0.984, 0.979, 0.974, 0.968, 0.962, 0.956, 
    0.95, 0.942, 0.935, 0.927, 0.918, 0.909, 0.899, 0.889, 0.879, 0.868, 
    0.857, 0.846, 0.835, 0.824, 0.814, 0.803, 0.793, 0.784, 0.774, 0.766, 
    0.757, 0.75, 0.743, 0.736, 0.73, 0.724, 0.719, 0.715, 0.711, 0.708, 
    0.705, 0.703, 0.701, 0.699, 0.699, 0.698, 0.699, 0.699, 0.7, 0.702, 
    0.704, 0.706, 0.709, 0.712, 0.715, 0.718, 0.722, 0.725, 0.729, 0.732, 
    0.736, 0.739, 0.743, 0.746, 0.749, 0.753, 0.757, 0.76, 0.764, 0.769, 
    0.774, 0.779, 0.785, 0.792, 0.799, 0.807, 0.816, 0.826, 0.837, 0.848, 
    0.86, 0.874, 0.888, 0.903, 0.919, 0.936, 0.954, 0.973, 0.994, 1.015, 
    1.038, 1.062, 1.088, 1.115, 1.145, 1.176, 1.209, 1.244, 1.282, 1.322, 
    1.364, 1.41, 1.458, 1.509, 1.564, 1.622, 1.683, 1.747, 1.815, 1.886, 
    1.96, 2.037, 2.116, 2.198, 2.28, 2.363, 2.445, 2.524, 2.601, 2.674, 
    2.741, 2.8, 2.851, 2.893, 2.925, 2.947, 2.959, 2.961, 2.954, 2.938, 
    2.916, 2.887, 2.853, 2.815, 2.773, 2.729, 2.683, 2.636, 2.587, 2.537, 
    2.484, 2.43, 2.377, 2.323, 2.272, 2.222, 2.177, 2.134, 2.092, 2.054, 
    2.017, 1.982, 1.947, 1.911, 1.875, 1.837, 1.801, 1.76, 1.716, 1.671, 
    1.621, 1.573, 1.521, 1.468, 1.417, 1.37, 1.328, 1.293, 1.267, 1.248, 
    1.235, 1.231, 1.238, 1.255, 1.281, 1.316, 1.36, 1.414, 1.477, 1.55, 
    1.632, 1.722, 1.819, 1.924, 2.038, 2.158, 2.284, 2.412, 2.536, 2.649, 
    2.738, 2.802, 2.839, 2.847, 2.83, 2.797, 2.751, 2.706, 2.657, 2.611, 
    2.562, 2.515, 2.465, 2.419, 2.371, 2.321, 2.273, 2.225, 2.179, 2.135, 
    2.092, 2.053, 2.014, 1.98, 1.951, 1.928, 1.914, 1.908, 1.913, 1.931, 
    1.962, 2.006, 2.063, 2.131, 2.204, 2.279, 2.351, 2.414, 2.464, 2.501, 
    2.528, 2.547, 2.559, 2.569, 2.577, 2.583, 2.591, 2.598, 2.603, 2.605, 
    2.604, 2.601, 2.596, 2.594, 2.594, 2.598, 2.606, 2.616, 2.626, 2.633, 
    2.633, 2.625, 2.608, 2.584, 2.556, 2.527, 2.498, 2.47, 2.443, 2.417, 
    2.393, 2.369, 2.347, 2.324, 2.301, 2.278, 2.258, 2.238, 2.219, 2.202, 
    2.184, 2.168, 2.153, 2.137, 2.123, 2.109, 2.096, 2.083, 2.072, 2.06, 
    2.049, 2.039, 2.03, 2.021, 2.013, 2.006, 2.001, 1.996, 1.993, 1.989, 
    1.985, 1.981, 1.972, 1.961, 1.944, 1.922, 1.897, 1.866, 1.833, 1.801, 
    1.766, 1.738, 1.719, 1.713, 1.724, 1.754, 1.804, 1.875, 1.965, 2.065, 
    2.167, 2.257, 2.323, 2.367, 2.391, 2.405, 2.415, 2.429, 2.447, 2.469, 
    2.493, 2.515, 2.534, 2.544, 2.549, 2.549, 2.542, 2.53, 2.516, 2.502, 
    2.491, 2.482, 2.476, 2.47, 2.466, 2.462, 2.459, 2.453, 2.444, 2.43, 
    2.414, 2.396, 2.378, 2.359, 2.341, 2.324, 2.308, 2.294, 2.282, 2.27, 
    2.26, 2.251, 2.24, 2.231, 2.221, 2.21, 2.197, 2.184, 2.17, 2.156, 2.141, 
    2.125, 2.11, 2.093, 2.075, 2.054, 2.033, 2.015, 1.998, 1.987, 1.977, 
    1.972, 1.975, 1.989, 2.014, 2.052, 2.102, 2.164, 2.238, 2.319, 2.401, 
    2.477, 2.538, 2.585, 2.618, 2.641, 2.656, 2.667, 2.674, 2.681, 2.683, 
    2.679, 2.669, 2.653, 2.632, 2.609, 2.585, 2.563, 2.542, 2.522, 2.503, 
    2.486, 2.469, 2.452, 2.438, 2.423, 2.411, 2.401, 2.392, 2.387, 2.383, 
    2.379, 2.375, 2.373, 2.37, 2.368, 2.367, 2.364, 2.363, 2.36, 2.357, 
    2.354, 2.351, 2.348, 2.345, 2.343, 2.339, 2.337, 2.335, 2.331, 2.328, 
    2.323, 2.319, 2.314, 2.307, 2.301, 2.295, 2.289, 2.283, 2.276, 2.268, 
    2.259, 2.249, 2.237, 2.226, 2.212, 2.199, 2.185, 2.172, 2.156, 2.139, 
    2.123, 2.108, 2.094, 2.083, 2.077, 2.076, 2.084, 2.102, 2.129, 2.164, 
    2.202, 2.241, 2.28, 2.313, 2.339, 2.358, 2.367, 2.372, 2.374, 2.376, 
    2.379, 2.38, 2.38, 2.381, 2.382, 2.382, 2.383, 2.382, 2.382, 2.382, 
    2.381, 2.38, 2.377, 2.373, 2.368, 2.362, 2.357, 2.351, 2.345, 2.339, 
    2.334, 2.328, 2.324, 2.319, 2.315, 2.311, 2.307, 2.304, 2.302, 2.299, 
    2.297, 2.295, 2.292, 2.289, 2.286, 2.283, 2.281, 2.279, 2.278, 2.278, 
    2.279, 2.281, 2.283, 2.285, 2.286, 2.287, 2.289, 2.29, 2.291, 2.293, 
    2.295, 2.296, 2.298, 2.302, 2.304, 2.308, 2.313, 2.319, 2.326, 2.333, 
    2.34, 2.349, 2.356, 2.364, 2.372, 2.382, 2.389, 2.395, 2.4, 2.404, 2.404, 
    2.403, 2.402, 2.4, 2.396, 2.392, 2.39, 2.387, 2.384, 2.38, 2.377, 2.373, 
    2.369, 2.365, 2.362, 2.358, 2.354, 2.349, 2.345, 2.341, 2.337, 2.333, 
    2.329, 2.324, 2.32, 2.316, 2.313, 2.31, 2.306, 2.303, 2.3, 2.296, 2.293, 
    2.289, 2.286, 2.282, 2.278, 2.275, 2.272, 2.269, 2.266, 2.263, 2.26, 
    2.256, 2.253, 2.249, 2.246, 2.246, 2.244, 2.244, 2.244, 2.245, 2.247, 
    2.25, 2.253, 2.257, 2.26, 2.264, 2.268, 2.272, 2.274, 2.277, 2.281, 
    2.284, 2.287 ;

 idx_rfr_kaolinite_img = 0.0009549926, 0.0001047129, 0.001202264, 
    0.001412538, 0.001258925, 0.001380385, 0.001230269, 0.001202264, 
    0.001230269, 0.001174897, 0.001174897, 0.001071519, 0.0008128307, 
    0.0003981071, 0.0002754229, 0.0002041738, 0.000144544, 0.0001230269, 
    9.549926e-05, 5.248072e-05, 3.890453e-05, 3.801893e-05, 4.168693e-05, 
    9.332538e-05, 1e-04, 0.0001288249, 0.0001230269, 0.0001584893, 
    0.0001348963, 0.0001584893, 0.0002041738, 0.0003467368, 0.0003090295, 
    0.0003162278, 0.0004073802, 0.0004570883, 0.0005623413, 0.0005623413, 
    0.0006918308, 0.001202264, 0.001778279, 0.001584893, 0.003311311, 
// NB: Relabel EgH79 value at 2.5 um as 2.4999 um to make room for 2.5 um Roush datum
// NB: Excise EgH79 value at 2.6 um in favor of Roush data
// end EgH79 Kaolinite. Begin Roush Kaolinite:
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001, 
    0.001, 0.002, 0.002, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.002, 
    0.002, 0.002, 0.001, 0.001, 0.001, 0.001, 0.002, 0.002, 0.002, 0.003, 
    0.004, 0.004, 0.004, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 
    0.005, 0.005, 0.005, 0.004, 0.004, 0.005, 0.004, 0.004, 0.004, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.004, 0.004, 0.005, 0.005, 
    0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.005, 0.005, 0.005, 
    0.004, 0.004, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.004, 
    0.004, 0.005, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 
    0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 
    0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 
    0.005, 0.006, 0.006, 0.007, 0.007, 0.008, 0.008, 0.009, 0.009, 0.009, 
    0.009, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.009, 0.009, 
    0.009, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.011, 0.011, 0.011, 0.011, 0.011, 0.01, 0.01, 
    0.009, 0.009, 0.008, 0.007, 0.007, 0.007, 0.007, 0.007, 0.008, 0.008, 
    0.009, 0.01, 0.01, 0.011, 0.011, 0.012, 0.012, 0.012, 0.011, 0.011, 
    0.011, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.011, 0.011, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.011, 0.011, 0.01, 0.01, 0.009, 
    0.009, 0.008, 0.008, 0.008, 0.008, 0.008, 0.007, 0.008, 0.007, 0.007, 
    0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.008, 0.008, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.011, 0.011, 0.011, 0.011, 0.011, 0.01, 
    0.01, 0.009, 0.008, 0.008, 0.007, 0.006, 0.006, 0.005, 0.005, 0.005, 
    0.005, 0.006, 0.006, 0.007, 0.008, 0.009, 0.01, 0.011, 0.012, 0.012, 
    0.012, 0.012, 0.011, 0.01, 0.01, 0.009, 0.009, 0.008, 0.008, 0.008, 
    0.008, 0.009, 0.01, 0.011, 0.012, 0.013, 0.015, 0.017, 0.019, 0.021, 
    0.023, 0.026, 0.029, 0.032, 0.035, 0.039, 0.042, 0.046, 0.049, 0.052, 
    0.056, 0.059, 0.061, 0.064, 0.065, 0.067, 0.067, 0.067, 0.067, 0.067, 
    0.066, 0.065, 0.065, 0.063, 0.063, 0.062, 0.061, 0.06, 0.059, 0.058, 
    0.057, 0.057, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.057, 
    0.058, 0.058, 0.059, 0.059, 0.06, 0.06, 0.06, 0.061, 0.061, 0.061, 0.061, 
    0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.06, 
    0.06, 0.06, 0.06, 0.059, 0.059, 0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 
    0.059, 0.06, 0.061, 0.064, 0.067, 0.071, 0.077, 0.083, 0.09, 0.098, 
    0.105, 0.112, 0.117, 0.122, 0.124, 0.125, 0.123, 0.119, 0.112, 0.105, 
    0.096, 0.086, 0.077, 0.068, 0.06, 0.053, 0.048, 0.044, 0.041, 0.04, 
    0.039, 0.038, 0.039, 0.039, 0.039, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.039, 0.039, 0.038, 0.037, 0.036, 0.035, 0.034, 0.034, 0.033, 0.033, 
    0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.033, 0.033, 0.033, 0.033, 
    0.033, 0.033, 0.033, 0.033, 0.033, 0.032, 0.032, 0.032, 0.033, 0.033, 
    0.033, 0.033, 0.033, 0.034, 0.034, 0.034, 0.035, 0.035, 0.035, 0.035, 
    0.036, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.034, 0.034, 0.034, 
    0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.034, 
    0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.033, 0.033, 
    0.033, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 
    0.033, 0.033, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.033, 
    0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 
    0.033, 0.033, 0.033, 0.033, 0.034, 0.034, 0.034, 0.034, 0.034, 0.035, 
    0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.036, 
    0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 
    0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 
    0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 
    0.036, 0.036, 0.036, 0.036, 0.036, 0.037, 0.037, 0.037, 0.037, 0.037, 
    0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 
    0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 
    0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 
    0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 
    0.037, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.04, 0.04, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.043, 0.043, 0.043, 0.043, 0.042, 0.042, 
    0.042, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.048, 
    0.048, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 
    0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 
    0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 
    0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.052, 0.052, 0.052, 0.052, 
    0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 
    0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 
    0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 
    0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 
    0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.056, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.054, 0.054, 0.054, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.054, 0.054, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.054, 0.054, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.054, 0.054, 0.054, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.054, 0.054, 0.054, 0.054, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.054, 0.054, 0.054, 0.054, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.054, 0.054, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.054, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 
    0.055, 0.055, 0.055, 0.055, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 
    0.056, 0.055, 0.055, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 
    0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 
    0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 
    0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 
    0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 
    0.056, 0.056, 0.056, 0.056, 0.056, 0.057, 0.057, 0.057, 0.057, 0.057, 
    0.057, 0.056, 0.056, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 
    0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 
    0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 
    0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 
    0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.058, 0.058, 0.058, 
    0.058, 0.057, 0.057, 0.058, 0.058, 0.058, 0.057, 0.057, 0.058, 0.058, 
    0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 
    0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 0.059, 0.059, 
    0.059, 0.058, 0.058, 0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 
    0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 
    0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.06, 0.06, 0.06, 
    0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 
    0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 0.061, 
    0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 
    0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.062, 0.062, 0.062, 0.062, 
    0.062, 0.062, 0.062, 0.062, 0.062, 0.062, 0.062, 0.062, 0.062, 0.062, 
    0.062, 0.062, 0.063, 0.063, 0.063, 0.063, 0.063, 0.062, 0.062, 0.063, 
    0.063, 0.063, 0.063, 0.063, 0.063, 0.063, 0.063, 0.063, 0.063, 0.063, 
    0.063, 0.063, 0.064, 0.064, 0.064, 0.064, 0.064, 0.064, 0.064, 0.064, 
    0.064, 0.064, 0.064, 0.064, 0.064, 0.064, 0.064, 0.064, 0.064, 0.065, 
    0.065, 0.065, 0.065, 0.065, 0.065, 0.065, 0.065, 0.065, 0.065, 0.065, 
    0.065, 0.065, 0.065, 0.065, 0.065, 0.065, 0.065, 0.065, 0.065, 0.065, 
    0.065, 0.065, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 
    0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 
    0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 
    0.067, 0.067, 0.067, 0.067, 0.066, 0.066, 0.066, 0.066, 0.066, 0.067, 
    0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.066, 0.066, 0.067, 0.067, 
    0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 
    0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 
    0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 
    0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 
    0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 
    0.067, 0.067, 0.067, 0.067, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.067, 0.067, 0.068, 0.068, 0.068, 0.067, 0.067, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.067, 0.068, 0.068, 
    0.068, 0.067, 0.068, 0.067, 0.067, 0.067, 0.067, 0.067, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.067, 0.068, 0.067, 0.067, 0.068, 0.067, 0.067, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.067, 0.068, 0.068, 0.067, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.068, 0.068, 0.069, 0.069, 0.068, 0.069, 0.069, 
    0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 
    0.069, 0.07, 0.069, 0.069, 0.07, 0.069, 0.069, 0.07, 0.07, 0.07, 0.07, 
    0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 
    0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 
    0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 
    0.07, 0.07, 0.07, 0.071, 0.07, 0.07, 0.07, 0.07, 0.071, 0.07, 0.07, 
    0.071, 0.07, 0.071, 0.071, 0.07, 0.071, 0.07, 0.07, 0.07, 0.07, 0.07, 
    0.071, 0.07, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 
    0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 
    0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 
    0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 
    0.071, 0.071, 0.071, 0.071, 0.072, 0.071, 0.072, 0.072, 0.072, 0.072, 
    0.072, 0.072, 0.072, 0.071, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 
    0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 
    0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 
    0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.071, 0.071, 0.072, 0.072, 
    0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 
    0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 
    0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 
    0.072, 0.072, 0.072, 0.072, 0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 
    0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 
    0.073, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 
    0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.075, 0.074, 
    0.074, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.076, 0.076, 0.076, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.076, 0.076, 0.076, 0.076, 0.076, 0.076, 0.076, 
    0.076, 0.076, 0.076, 0.076, 0.076, 0.076, 0.076, 0.076, 0.076, 0.076, 
    0.076, 0.077, 0.077, 0.077, 0.077, 0.077, 0.077, 0.077, 0.077, 0.078, 
    0.078, 0.077, 0.077, 0.077, 0.077, 0.077, 0.077, 0.077, 0.077, 0.077, 
    0.077, 0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 
    0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 
    0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 0.078, 
    0.078, 0.077, 0.077, 0.078, 0.077, 0.078, 0.078, 0.078, 0.079, 0.079, 
    0.08, 0.08, 0.08, 0.081, 0.081, 0.082, 0.082, 0.082, 0.083, 0.083, 0.083, 
    0.084, 0.085, 0.085, 0.085, 0.085, 0.086, 0.086, 0.086, 0.087, 0.087, 
    0.087, 0.087, 0.087, 0.088, 0.088, 0.088, 0.088, 0.088, 0.088, 0.088, 
    0.087, 0.087, 0.087, 0.087, 0.087, 0.087, 0.087, 0.088, 0.087, 0.087, 
    0.088, 0.088, 0.088, 0.088, 0.088, 0.088, 0.088, 0.088, 0.088, 0.088, 
    0.088, 0.088, 0.088, 0.088, 0.088, 0.088, 0.088, 0.088, 0.088, 0.088, 
    0.088, 0.089, 0.089, 0.089, 0.09, 0.09, 0.09, 0.091, 0.091, 0.091, 0.092, 
    0.092, 0.092, 0.092, 0.092, 0.092, 0.093, 0.093, 0.093, 0.093, 0.094, 
    0.094, 0.094, 0.094, 0.095, 0.095, 0.095, 0.096, 0.096, 0.096, 0.096, 
    0.096, 0.096, 0.096, 0.096, 0.097, 0.097, 0.097, 0.097, 0.097, 0.097, 
    0.097, 0.097, 0.097, 0.097, 0.098, 0.097, 0.098, 0.099, 0.099, 0.1, 
    0.101, 0.102, 0.102, 0.103, 0.104, 0.105, 0.106, 0.106, 0.107, 0.107, 
    0.107, 0.108, 0.109, 0.109, 0.11, 0.11, 0.11, 0.111, 0.111, 0.111, 0.111, 
    0.111, 0.112, 0.112, 0.112, 0.113, 0.113, 0.114, 0.114, 0.115, 0.116, 
    0.117, 0.117, 0.118, 0.118, 0.119, 0.12, 0.121, 0.122, 0.123, 0.124, 
    0.125, 0.126, 0.127, 0.128, 0.13, 0.131, 0.132, 0.134, 0.135, 0.137, 
    0.138, 0.139, 0.141, 0.142, 0.143, 0.144, 0.145, 0.146, 0.148, 0.149, 
    0.15, 0.152, 0.154, 0.156, 0.159, 0.162, 0.166, 0.171, 0.177, 0.183, 
    0.191, 0.199, 0.208, 0.218, 0.23, 0.242, 0.255, 0.268, 0.283, 0.299, 
    0.315, 0.332, 0.35, 0.369, 0.388, 0.408, 0.429, 0.45, 0.471, 0.493, 
    0.515, 0.537, 0.558, 0.579, 0.6, 0.62, 0.638, 0.655, 0.671, 0.684, 0.695, 
    0.702, 0.707, 0.709, 0.707, 0.702, 0.694, 0.683, 0.67, 0.656, 0.64, 
    0.623, 0.607, 0.592, 0.578, 0.566, 0.556, 0.548, 0.543, 0.54, 0.54, 
    0.543, 0.547, 0.554, 0.563, 0.575, 0.588, 0.603, 0.619, 0.637, 0.657, 
    0.677, 0.699, 0.722, 0.746, 0.771, 0.797, 0.823, 0.851, 0.878, 0.906, 
    0.935, 0.964, 0.993, 1.02, 1.05, 1.08, 1.11, 1.14, 1.17, 1.2, 1.23, 1.26, 
    1.29, 1.32, 1.36, 1.39, 1.42, 1.45, 1.48, 1.51, 1.55, 1.58, 1.61, 1.65, 
    1.68, 1.72, 1.75, 1.79, 1.83, 1.87, 1.91, 1.95, 1.99, 2.03, 2.07, 2.12, 
    2.16, 2.2, 2.24, 2.27, 2.3, 2.33, 2.35, 2.36, 2.35, 2.34, 2.32, 2.28, 
    2.24, 2.18, 2.12, 2.05, 1.98, 1.91, 1.85, 1.78, 1.72, 1.66, 1.61, 1.56, 
    1.52, 1.48, 1.45, 1.42, 1.4, 1.37, 1.36, 1.34, 1.33, 1.31, 1.3, 1.29, 
    1.28, 1.27, 1.25, 1.24, 1.22, 1.19, 1.16, 1.13, 1.09, 1.03, 0.978, 0.914, 
    0.845, 0.77, 0.695, 0.618, 0.543, 0.472, 0.407, 0.347, 0.296, 0.252, 
    0.216, 0.187, 0.164, 0.147, 0.135, 0.126, 0.121, 0.118, 0.117, 0.116, 
    0.117, 0.119, 0.12, 0.122, 0.124, 0.127, 0.129, 0.132, 0.135, 0.139, 
    0.144, 0.149, 0.155, 0.162, 0.17, 0.179, 0.189, 0.199, 0.211, 0.223, 
    0.236, 0.25, 0.264, 0.278, 0.292, 0.307, 0.321, 0.335, 0.349, 0.363, 
    0.377, 0.391, 0.404, 0.418, 0.431, 0.444, 0.458, 0.471, 0.485, 0.5, 
    0.515, 0.53, 0.545, 0.561, 0.578, 0.594, 0.611, 0.628, 0.644, 0.66, 
    0.676, 0.69, 0.704, 0.717, 0.728, 0.738, 0.746, 0.753, 0.758, 0.761, 
    0.762, 0.761, 0.757, 0.751, 0.743, 0.732, 0.718, 0.701, 0.682, 0.659, 
    0.633, 0.605, 0.574, 0.541, 0.506, 0.47, 0.434, 0.398, 0.363, 0.329, 
    0.297, 0.267, 0.24, 0.215, 0.194, 0.175, 0.159, 0.146, 0.135, 0.126, 
    0.119, 0.113, 0.109, 0.105, 0.102, 0.1, 0.098, 0.096, 0.094, 0.092, 0.09, 
    0.088, 0.086, 0.084, 0.082, 0.081, 0.079, 0.077, 0.076, 0.075, 0.073, 
    0.072, 0.071, 0.07, 0.069, 0.068, 0.067, 0.067, 0.066, 0.065, 0.065, 
    0.064, 0.064, 0.063, 0.063, 0.063, 0.063, 0.062, 0.062, 0.062, 0.062, 
    0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 
    0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.061, 0.062, 0.062, 0.062, 
    0.062, 0.063, 0.064, 0.064, 0.065, 0.066, 0.068, 0.069, 0.071, 0.074, 
    0.077, 0.08, 0.083, 0.087, 0.091, 0.095, 0.099, 0.104, 0.109, 0.113, 
    0.119, 0.124, 0.128, 0.133, 0.138, 0.143, 0.147, 0.151, 0.155, 0.159, 
    0.162, 0.165, 0.167, 0.169, 0.171, 0.172, 0.173, 0.173, 0.172, 0.172, 
    0.17, 0.168, 0.166, 0.164, 0.161, 0.158, 0.154, 0.151, 0.148, 0.144, 
    0.141, 0.138, 0.136, 0.133, 0.131, 0.13, 0.128, 0.127, 0.127, 0.127, 
    0.127, 0.128, 0.129, 0.13, 0.132, 0.133, 0.135, 0.137, 0.14, 0.142, 
    0.144, 0.146, 0.147, 0.149, 0.151, 0.152, 0.153, 0.154, 0.155, 0.155, 
    0.156, 0.156, 0.156, 0.155, 0.155, 0.154, 0.153, 0.151, 0.15, 0.148, 
    0.146, 0.144, 0.142, 0.139, 0.137, 0.135, 0.133, 0.131, 0.129, 0.127, 
    0.126, 0.125, 0.124, 0.123, 0.123, 0.124, 0.124, 0.126, 0.127, 0.13, 
    0.132, 0.135, 0.138, 0.142, 0.146, 0.15, 0.154, 0.159, 0.164, 0.168, 
    0.174, 0.178, 0.184, 0.189, 0.195, 0.2, 0.206, 0.211, 0.217, 0.222, 
    0.227, 0.232, 0.237, 0.242, 0.247, 0.251, 0.255, 0.259, 0.263, 0.266, 
    0.27, 0.272, 0.275, 0.277, 0.28, 0.282, 0.284, 0.286, 0.287, 0.289, 0.29, 
    0.292, 0.294, 0.295, 0.297, 0.299, 0.301, 0.303, 0.305, 0.307, 0.31, 
    0.313, 0.316, 0.32, 0.323, 0.327, 0.33, 0.335, 0.339, 0.343, 0.347, 
    0.352, 0.356, 0.36, 0.364, 0.368, 0.371, 0.375, 0.379, 0.382, 0.385, 
    0.388, 0.391, 0.394, 0.398, 0.401, 0.404, 0.408, 0.412, 0.417, 0.422, 
    0.428, 0.434, 0.441, 0.449, 0.458, 0.467, 0.478, 0.489, 0.501, 0.514, 
    0.527, 0.541, 0.556, 0.571, 0.587, 0.603, 0.619, 0.636, 0.653, 0.67, 
    0.688, 0.706, 0.724, 0.742, 0.76, 0.778, 0.797, 0.815, 0.834, 0.852, 
    0.87, 0.889, 0.907, 0.925, 0.943, 0.961, 0.979, 0.996, 1.01, 1.03, 1.05, 
    1.07, 1.08, 1.1, 1.12, 1.13, 1.15, 1.17, 1.19, 1.21, 1.23, 1.25, 1.27, 
    1.29, 1.31, 1.33, 1.36, 1.38, 1.4, 1.43, 1.45, 1.48, 1.5, 1.53, 1.55, 
    1.58, 1.61, 1.63, 1.66, 1.69, 1.71, 1.74, 1.77, 1.79, 1.82, 1.85, 1.88, 
    1.91, 1.94, 1.96, 1.99, 2.02, 2.05, 2.07, 2.1, 2.12, 2.15, 2.17, 2.19, 
    2.21, 2.22, 2.23, 2.24, 2.24, 2.24, 2.23, 2.21, 2.19, 2.16, 2.12, 2.07, 
    2.02, 1.95, 1.88, 1.8, 1.72, 1.63, 1.53, 1.44, 1.35, 1.25, 1.16, 1.07, 
    0.991, 0.913, 0.842, 0.776, 0.716, 0.661, 0.611, 0.566, 0.525, 0.489, 
    0.456, 0.43, 0.409, 0.393, 0.383, 0.377, 0.375, 0.374, 0.375, 0.378, 
    0.381, 0.383, 0.385, 0.388, 0.391, 0.396, 0.401, 0.405, 0.413, 0.424, 
    0.439, 0.461, 0.485, 0.519, 0.562, 0.613, 0.672, 0.74, 0.812, 0.886, 
    0.965, 1.05, 1.13, 1.22, 1.3, 1.38, 1.46, 1.53, 1.6, 1.67, 1.73, 1.77, 
    1.81, 1.85, 1.86, 1.87, 1.85, 1.82, 1.75, 1.66, 1.55, 1.43, 1.3, 1.17, 
    1.06, 0.957, 0.877, 0.811, 0.756, 0.711, 0.671, 0.64, 0.613, 0.594, 
    0.576, 0.566, 0.562, 0.564, 0.571, 0.583, 0.601, 0.624, 0.652, 0.687, 
    0.729, 0.777, 0.829, 0.887, 0.949, 1.01, 1.07, 1.13, 1.17, 1.21, 1.23, 
    1.23, 1.21, 1.18, 1.14, 1.1, 1.05, 1.01, 0.974, 0.941, 0.911, 0.883, 
    0.857, 0.83, 0.802, 0.773, 0.747, 0.723, 0.702, 0.686, 0.67, 0.654, 
    0.637, 0.615, 0.587, 0.553, 0.513, 0.472, 0.431, 0.396, 0.367, 0.344, 
    0.326, 0.312, 0.3, 0.292, 0.285, 0.279, 0.274, 0.27, 0.268, 0.269, 0.27, 
    0.272, 0.276, 0.279, 0.283, 0.289, 0.294, 0.299, 0.306, 0.313, 0.321, 
    0.328, 0.337, 0.345, 0.354, 0.364, 0.373, 0.383, 0.393, 0.403, 0.414, 
    0.422, 0.431, 0.437, 0.441, 0.444, 0.444, 0.444, 0.445, 0.447, 0.454, 
    0.467, 0.487, 0.516, 0.553, 0.606, 0.668, 0.743, 0.824, 0.908, 0.988, 
    1.06, 1.11, 1.13, 1.13, 1.1, 1.04, 0.992, 0.941, 0.903, 0.875, 0.856, 
    0.838, 0.82, 0.795, 0.766, 0.73, 0.693, 0.655, 0.619, 0.585, 0.555, 
    0.531, 0.513, 0.499, 0.488, 0.476, 0.464, 0.451, 0.437, 0.422, 0.404, 
    0.385, 0.366, 0.351, 0.339, 0.329, 0.322, 0.318, 0.316, 0.316, 0.317, 
    0.319, 0.32, 0.322, 0.324, 0.324, 0.325, 0.325, 0.325, 0.326, 0.328, 
    0.331, 0.334, 0.34, 0.347, 0.355, 0.364, 0.375, 0.39, 0.411, 0.437, 
    0.468, 0.503, 0.54, 0.586, 0.636, 0.69, 0.745, 0.799, 0.847, 0.887, 
    0.915, 0.926, 0.916, 0.888, 0.843, 0.792, 0.74, 0.689, 0.641, 0.597, 
    0.556, 0.515, 0.473, 0.43, 0.389, 0.352, 0.32, 0.294, 0.274, 0.258, 
    0.245, 0.236, 0.228, 0.222, 0.217, 0.214, 0.213, 0.214, 0.216, 0.219, 
    0.223, 0.227, 0.228, 0.229, 0.23, 0.231, 0.231, 0.23, 0.229, 0.227, 
    0.225, 0.222, 0.219, 0.217, 0.214, 0.211, 0.209, 0.206, 0.204, 0.201, 
    0.197, 0.193, 0.189, 0.185, 0.181, 0.177, 0.173, 0.171, 0.168, 0.165, 
    0.162, 0.158, 0.155, 0.152, 0.149, 0.148, 0.148, 0.148, 0.151, 0.156, 
    0.161, 0.166, 0.177, 0.191, 0.208, 0.23, 0.256, 0.286, 0.319, 0.355, 
    0.39, 0.421, 0.444, 0.458, 0.462, 0.458, 0.444, 0.424, 0.401, 0.378, 
    0.358, 0.342, 0.329, 0.318, 0.307, 0.297, 0.288, 0.279, 0.271, 0.262, 
    0.254, 0.246, 0.238, 0.23, 0.221, 0.211, 0.203, 0.196, 0.19, 0.184, 0.18, 
    0.176, 0.174, 0.172, 0.17, 0.169, 0.169, 0.168, 0.168, 0.168, 0.169, 
    0.17, 0.17, 0.17, 0.171, 0.171, 0.172, 0.173, 0.175, 0.177, 0.18, 0.184, 
    0.187, 0.191, 0.193, 0.195, 0.196, 0.197, 0.198, 0.199, 0.2, 0.201, 
    0.203, 0.204, 0.206, 0.208, 0.21, 0.212, 0.214, 0.217, 0.219, 0.219, 
    0.219, 0.219, 0.217, 0.214, 0.21, 0.206, 0.2, 0.191, 0.182, 0.171, 0.16, 
    0.148, 0.138, 0.129, 0.12, 0.111, 0.105, 0.099, 0.093, 0.087, 0.081, 
    0.076, 0.071, 0.067, 0.063, 0.059, 0.055, 0.051, 0.047, 0.045, 0.042, 
    0.04, 0.038, 0.036, 0.034, 0.033, 0.032, 0.031, 0.03, 0.029, 0.028, 
    0.028, 0.027, 0.026, 0.026, 0.026, 0.026, 0.026, 0.027, 0.028, 0.028, 
    0.029, 0.03, 0.031, 0.033, 0.035, 0.038, 0.042, 0.046, 0.05, 0.054, 
    0.059, 0.063, 0.067, 0.07, 0.073, 0.075, 0.076, 0.077, 0.077, 0.076, 
    0.075, 0.074, 0.073, 0.07, 0.067 ;

 bnd_montmorillonite = 0.185, 0.19, 0.2, 0.21, 0.215, 0.22, 0.225, 0.233, 0.24, 0.26, 0.28, 
    0.3, 0.325, 0.36, 0.37, 0.4, 0.433, 0.466, 0.5, 0.533, 0.566, 0.6, 0.633, 
    0.666, 0.7, 0.817, 0.907, 1, 1.105, 1.2, 1.303, 1.4, 1.5, 1.6, 1.7, 1.8, 
    1.9, 2, 2.1, 2.2, 2.3, 2.4, 2.4999,
    5, 5.01, 5.02, 5.03, 5.04, 5.05, 5.061, 5.071, 5.081, 5.092, 5.102, 
    5.113, 5.123, 5.134, 5.144, 5.155, 5.165, 5.176, 5.187, 5.198, 5.208, 
    5.219, 5.23, 5.241, 5.252, 5.263, 5.274, 5.285, 5.297, 5.308, 5.319, 
    5.331, 5.342, 5.353, 5.365, 5.376, 5.388, 5.4, 5.411, 5.423, 5.435, 
    5.447, 5.458, 5.47, 5.483, 5.495, 5.507, 5.519, 5.531, 5.543, 5.556, 
    5.568, 5.58, 5.593, 5.605, 5.618, 5.631, 5.643, 5.656, 5.669, 5.682, 
    5.695, 5.708, 5.721, 5.734, 5.747, 5.76, 5.774, 5.787, 5.8, 5.814, 5.827, 
    5.841, 5.855, 5.869, 5.882, 5.896, 5.91, 5.924, 5.938, 5.952, 5.967, 
    5.981, 5.995, 6.01, 6.024, 6.039, 6.053, 6.068, 6.083, 6.098, 6.113, 
    6.128, 6.142, 6.158, 6.173, 6.188, 6.203, 6.219, 6.234, 6.25, 6.266, 
    6.281, 6.297, 6.313, 6.329, 6.345, 6.361, 6.378, 6.394, 6.41, 6.427, 
    6.443, 6.46, 6.477, 6.494, 6.51, 6.527, 6.544, 6.562, 6.579, 6.596, 
    6.614, 6.631, 6.649, 6.667, 6.685, 6.702, 6.72, 6.739, 6.757, 6.775, 
    6.793, 6.812, 6.831, 6.849, 6.868, 6.887, 6.906, 6.925, 6.944, 6.964, 
    6.983, 7.003, 7.023, 7.042, 7.062, 7.082, 7.102, 7.122, 7.143, 7.163, 
    7.184, 7.205, 7.225, 7.246, 7.267, 7.289, 7.31, 7.331, 7.353, 7.375, 
    7.396, 7.418, 7.44, 7.463, 7.485, 7.508, 7.53, 7.553, 7.576, 7.599, 
    7.622, 7.645, 7.669, 7.692, 7.716, 7.74, 7.764, 7.788, 7.813, 7.837, 
    7.862, 7.886, 7.911, 7.937, 7.962, 7.987, 8.013, 8.039, 8.064, 8.091, 
    8.117, 8.143, 8.17, 8.197, 8.224, 8.251, 8.278, 8.306, 8.333, 8.361, 
    8.389, 8.417, 8.446, 8.475, 8.503, 8.532, 8.562, 8.591, 8.621, 8.651, 
    8.681, 8.711, 8.741, 8.772, 8.803, 8.834, 8.865, 8.897, 8.929, 8.961, 
    8.993, 9.025, 9.058, 9.091, 9.124, 9.158, 9.191, 9.225, 9.259, 9.294, 
    9.328, 9.363, 9.399, 9.434, 9.47, 9.506, 9.542, 9.578, 9.615, 9.653, 
    9.69, 9.728, 9.766, 9.804, 9.842, 9.881, 9.921, 9.96, 10, 10.04, 10.081, 
    10.121, 10.163, 10.204, 10.246, 10.288, 10.331, 10.373, 10.417, 10.46, 
    10.504, 10.549, 10.593, 10.638, 10.684, 10.73, 10.776, 10.823, 10.87, 
    10.917, 10.965, 11.013, 11.062, 11.111, 11.161, 11.211, 11.261, 11.312, 
    11.364, 11.416, 11.468, 11.521, 11.574, 11.628, 11.682, 11.737, 11.792, 
    11.848, 11.905, 11.962, 12.019, 12.077, 12.136, 12.195, 12.255, 12.315, 
    12.376, 12.438, 12.5, 12.563, 12.626, 12.69, 12.755, 12.821, 12.887, 
    12.953, 13.021, 13.089, 13.158, 13.228, 13.298, 13.369, 13.441, 13.514, 
    13.587, 13.661, 13.736, 13.812, 13.889, 13.966, 14.045, 14.124, 14.205, 
    14.286, 14.368, 14.451, 14.535, 14.62, 14.706, 14.793, 14.881, 14.97, 
    15.06, 15.152, 15.244, 15.337, 15.432, 15.528, 15.625, 15.723, 15.823, 
    15.924, 16.026, 16.129, 16.234, 16.34, 16.447, 16.556, 16.667, 16.779, 
    16.892, 17.007, 17.123, 17.241, 17.361, 17.483, 17.606, 17.731, 17.857, 
    17.986, 18.116, 18.248, 18.382, 18.519, 18.657, 18.797, 18.939, 19.084, 
    19.231, 19.38, 19.531, 19.685, 19.841, 20, 20.161, 20.325, 20.492, 
    20.661, 20.833, 21.008, 21.186, 21.368, 21.552, 21.739, 21.93, 22.124, 
    22.321, 22.523, 22.727, 22.936, 23.148, 23.364, 23.585, 23.81, 24.038, 
    24.272, 24.51, 24.752, 25 ;

 idx_rfr_montmorillonite_rl = 1.544, 1.543, 1.542, 1.541, 1.54, 1.539, 1.539, 
    1.538, 1.537, 1.536, 1.534, 1.523, 1.523, 1.524, 1.524, 1.525, 1.525, 
    1.526, 1.526, 1.524, 1.522, 1.52, 1.522, 1.523, 1.525, 1.527, 1.528, 
    1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 
    1.53, 1.53, 1.53, 1.53,
    1.336, 1.335, 1.335, 1.335, 1.334, 1.334, 
    1.333, 1.333, 1.333, 1.332, 1.332, 1.332, 1.331, 1.331, 1.33, 1.33, 
    1.329, 1.329, 1.329, 1.328, 1.328, 1.327, 1.327, 1.326, 1.326, 1.325, 
    1.325, 1.324, 1.324, 1.324, 1.323, 1.322, 1.322, 1.321, 1.321, 1.32, 
    1.32, 1.319, 1.319, 1.318, 1.318, 1.317, 1.317, 1.316, 1.316, 1.315, 
    1.314, 1.314, 1.313, 1.313, 1.312, 1.311, 1.311, 1.31, 1.309, 1.309, 
    1.308, 1.308, 1.307, 1.306, 1.305, 1.305, 1.304, 1.303, 1.302, 1.302, 
    1.301, 1.3, 1.299, 1.298, 1.298, 1.297, 1.296, 1.295, 1.294, 1.293, 
    1.292, 1.291, 1.29, 1.289, 1.288, 1.287, 1.285, 1.284, 1.282, 1.281, 
    1.279, 1.276, 1.274, 1.271, 1.269, 1.272, 1.284, 1.294, 1.294, 1.291, 
    1.288, 1.286, 1.283, 1.281, 1.28, 1.278, 1.276, 1.275, 1.273, 1.271, 
    1.27, 1.269, 1.267, 1.266, 1.264, 1.263, 1.261, 1.26, 1.258, 1.257, 
    1.256, 1.254, 1.253, 1.251, 1.25, 1.248, 1.246, 1.245, 1.243, 1.241, 
    1.24, 1.238, 1.236, 1.234, 1.232, 1.231, 1.229, 1.227, 1.225, 1.223, 
    1.221, 1.219, 1.217, 1.214, 1.212, 1.21, 1.208, 1.205, 1.203, 1.201, 
    1.198, 1.195, 1.193, 1.19, 1.187, 1.185, 1.182, 1.179, 1.176, 1.173, 
    1.169, 1.166, 1.163, 1.159, 1.156, 1.152, 1.148, 1.145, 1.141, 1.137, 
    1.132, 1.128, 1.124, 1.119, 1.114, 1.109, 1.104, 1.099, 1.094, 1.088, 
    1.082, 1.076, 1.07, 1.063, 1.056, 1.049, 1.042, 1.034, 1.026, 1.018, 
    1.009, 1, 0.99, 0.98, 0.969, 0.957, 0.945, 0.933, 0.919, 0.905, 0.89, 
    0.874, 0.856, 0.838, 0.818, 0.797, 0.774, 0.75, 0.725, 0.699, 0.672, 
    0.645, 0.621, 0.6, 0.585, 0.577, 0.575, 0.579, 0.587, 0.601, 0.625, 
    0.663, 0.716, 0.777, 0.826, 0.844, 0.824, 0.779, 0.724, 0.671, 0.63, 
    0.605, 0.598, 0.609, 0.637, 0.684, 0.754, 0.851, 0.982, 1.153, 1.365, 
    1.601, 1.823, 1.986, 2.078, 2.126, 2.177, 2.259, 2.365, 2.458, 2.504, 
    2.501, 2.464, 2.409, 2.349, 2.289, 2.232, 2.179, 2.129, 2.084, 2.042, 
    2.003, 1.966, 1.932, 1.899, 1.868, 1.838, 1.809, 1.78, 1.752, 1.726, 
    1.706, 1.698, 1.713, 1.748, 1.777, 1.782, 1.769, 1.749, 1.727, 1.707, 
    1.692, 1.688, 1.695, 1.704, 1.705, 1.697, 1.682, 1.665, 1.648, 1.637, 
    1.642, 1.648, 1.639, 1.624, 1.61, 1.596, 1.583, 1.57, 1.558, 1.546, 
    1.533, 1.521, 1.51, 1.503, 1.505, 1.517, 1.527, 1.526, 1.518, 1.507, 
    1.495, 1.484, 1.474, 1.463, 1.453, 1.443, 1.433, 1.423, 1.412, 1.402, 
    1.392, 1.381, 1.37, 1.359, 1.347, 1.335, 1.323, 1.313, 1.308, 1.304, 
    1.294, 1.281, 1.266, 1.251, 1.235, 1.219, 1.203, 1.186, 1.169, 1.151, 
    1.133, 1.115, 1.097, 1.079, 1.062, 1.046, 1.031, 1.019, 1.009, 1.003, 
    0.999, 0.999, 1.001, 1.004, 1.007, 1.009, 1.008, 1.004, 0.999, 0.993, 
    0.992, 0.998, 1.018, 1.055, 1.109, 1.175, 1.247, 1.314, 1.383, 1.486, 
    1.674, 1.942, 2.143, 2.168, 2.08, 1.954, 1.817, 1.678, 1.538, 1.407, 
    1.315, 1.314, 1.451, 1.721, 2.019, 2.328, 2.744, 3.046, 3.073, 2.968, 
    2.843, 2.73, 2.634, 2.554, 2.486, 2.428, 2.379, 2.335, 2.297, 2.263, 
    2.233, 2.206, 2.181, 2.158 ;

 bnd_montmorillonite = 0.185, 0.19, 0.2, 0.21, 0.215, 0.22, 0.225, 0.233, 0.24, 0.26, 0.28, 
    0.3, 0.325, 0.36, 0.37, 0.4, 0.433, 0.466, 0.5, 0.533, 0.566, 0.6, 0.633, 
    0.666, 0.7, 0.817, 0.907, 1, 1.105, 1.2, 1.303, 1.4, 1.5, 1.6, 1.7, 1.8, 
    1.9, 2, 2.1, 2.2, 2.3, 2.4, 2.4999,
// NB: Relabel EgH79 value at 2.5 um as 2.4999 um to make room for 2.5 um Roush datum
// NB: Excise EgH79 value at 2.6 um in favor of Roush data
// end EgH79 Montmorillonite. Begin Roush Montmorillonite:
    5, 5.01, 5.02, 5.03, 5.04, 5.05, 5.061, 5.071, 5.081, 5.092, 5.102, 
    5.113, 5.123, 5.134, 5.144, 5.155, 5.165, 5.176, 5.187, 5.198, 5.208, 
    5.219, 5.23, 5.241, 5.252, 5.263, 5.274, 5.285, 5.297, 5.308, 5.319, 
    5.331, 5.342, 5.353, 5.365, 5.376, 5.388, 5.4, 5.411, 5.423, 5.435, 
    5.447, 5.458, 5.47, 5.483, 5.495, 5.507, 5.519, 5.531, 5.543, 5.556, 
    5.568, 5.58, 5.593, 5.605, 5.618, 5.631, 5.643, 5.656, 5.669, 5.682, 
    5.695, 5.708, 5.721, 5.734, 5.747, 5.76, 5.774, 5.787, 5.8, 5.814, 5.827, 
    5.841, 5.855, 5.869, 5.882, 5.896, 5.91, 5.924, 5.938, 5.952, 5.967, 
    5.981, 5.995, 6.01, 6.024, 6.039, 6.053, 6.068, 6.083, 6.098, 6.113, 
    6.128, 6.142, 6.158, 6.173, 6.188, 6.203, 6.219, 6.234, 6.25, 6.266, 
    6.281, 6.297, 6.313, 6.329, 6.345, 6.361, 6.378, 6.394, 6.41, 6.427, 
    6.443, 6.46, 6.477, 6.494, 6.51, 6.527, 6.544, 6.562, 6.579, 6.596, 
    6.614, 6.631, 6.649, 6.667, 6.685, 6.702, 6.72, 6.739, 6.757, 6.775, 
    6.793, 6.812, 6.831, 6.849, 6.868, 6.887, 6.906, 6.925, 6.944, 6.964, 
    6.983, 7.003, 7.023, 7.042, 7.062, 7.082, 7.102, 7.122, 7.143, 7.163, 
    7.184, 7.205, 7.225, 7.246, 7.267, 7.289, 7.31, 7.331, 7.353, 7.375, 
    7.396, 7.418, 7.44, 7.463, 7.485, 7.508, 7.53, 7.553, 7.576, 7.599, 
    7.622, 7.645, 7.669, 7.692, 7.716, 7.74, 7.764, 7.788, 7.813, 7.837, 
    7.862, 7.886, 7.911, 7.937, 7.962, 7.987, 8.013, 8.039, 8.064, 8.091, 
    8.117, 8.143, 8.17, 8.197, 8.224, 8.251, 8.278, 8.306, 8.333, 8.361, 
    8.389, 8.417, 8.446, 8.475, 8.503, 8.532, 8.562, 8.591, 8.621, 8.651, 
    8.681, 8.711, 8.741, 8.772, 8.803, 8.834, 8.865, 8.897, 8.929, 8.961, 
    8.993, 9.025, 9.058, 9.091, 9.124, 9.158, 9.191, 9.225, 9.259, 9.294, 
    9.328, 9.363, 9.399, 9.434, 9.47, 9.506, 9.542, 9.578, 9.615, 9.653, 
    9.69, 9.728, 9.766, 9.804, 9.842, 9.881, 9.921, 9.96, 10, 10.04, 10.081, 
    10.121, 10.163, 10.204, 10.246, 10.288, 10.331, 10.373, 10.417, 10.46, 
    10.504, 10.549, 10.593, 10.638, 10.684, 10.73, 10.776, 10.823, 10.87, 
    10.917, 10.965, 11.013, 11.062, 11.111, 11.161, 11.211, 11.261, 11.312, 
    11.364, 11.416, 11.468, 11.521, 11.574, 11.628, 11.682, 11.737, 11.792, 
    11.848, 11.905, 11.962, 12.019, 12.077, 12.136, 12.195, 12.255, 12.315, 
    12.376, 12.438, 12.5, 12.563, 12.626, 12.69, 12.755, 12.821, 12.887, 
    12.953, 13.021, 13.089, 13.158, 13.228, 13.298, 13.369, 13.441, 13.514, 
    13.587, 13.661, 13.736, 13.812, 13.889, 13.966, 14.045, 14.124, 14.205, 
    14.286, 14.368, 14.451, 14.535, 14.62, 14.706, 14.793, 14.881, 14.97, 
    15.06, 15.152, 15.244, 15.337, 15.432, 15.528, 15.625, 15.723, 15.823, 
    15.924, 16.026, 16.129, 16.234, 16.34, 16.447, 16.556, 16.667, 16.779, 
    16.892, 17.007, 17.123, 17.241, 17.361, 17.483, 17.606, 17.731, 17.857, 
    17.986, 18.116, 18.248, 18.382, 18.519, 18.657, 18.797, 18.939, 19.084, 
    19.231, 19.38, 19.531, 19.685, 19.841, 20, 20.161, 20.325, 20.492, 
    20.661, 20.833, 21.008, 21.186, 21.368, 21.552, 21.739, 21.93, 22.124, 
    22.321, 22.523, 22.727, 22.936, 23.148, 23.364, 23.585, 23.81, 24.038, 
    24.272, 24.51, 24.752, 25 ;

 idx_rfr_montmorillonite_rl = 1.544, 1.543, 1.542, 1.541, 1.54, 1.539, 1.539, 
    1.538, 1.537, 1.536, 1.534, 1.523, 1.523, 1.524, 1.524, 1.525, 1.525, 
    1.526, 1.526, 1.524, 1.522, 1.52, 1.522, 1.523, 1.525, 1.527, 1.528, 
    1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 
    1.53, 1.53, 1.53, 1.53,
// NB: Relabel EgH79 value at 2.5 um as 2.4999 um to make room for 2.5 um Roush datum
// NB: Excise EgH79 value at 2.6 um in favor of Roush data
// end EgH79 Montmorillonite. Begin Roush Montmorillonite:
    1.336, 1.335, 1.335, 1.335, 1.334, 1.334, 
    1.333, 1.333, 1.333, 1.332, 1.332, 1.332, 1.331, 1.331, 1.33, 1.33, 
    1.329, 1.329, 1.329, 1.328, 1.328, 1.327, 1.327, 1.326, 1.326, 1.325, 
    1.325, 1.324, 1.324, 1.324, 1.323, 1.322, 1.322, 1.321, 1.321, 1.32, 
    1.32, 1.319, 1.319, 1.318, 1.318, 1.317, 1.317, 1.316, 1.316, 1.315, 
    1.314, 1.314, 1.313, 1.313, 1.312, 1.311, 1.311, 1.31, 1.309, 1.309, 
    1.308, 1.308, 1.307, 1.306, 1.305, 1.305, 1.304, 1.303, 1.302, 1.302, 
    1.301, 1.3, 1.299, 1.298, 1.298, 1.297, 1.296, 1.295, 1.294, 1.293, 
    1.292, 1.291, 1.29, 1.289, 1.288, 1.287, 1.285, 1.284, 1.282, 1.281, 
    1.279, 1.276, 1.274, 1.271, 1.269, 1.272, 1.284, 1.294, 1.294, 1.291, 
    1.288, 1.286, 1.283, 1.281, 1.28, 1.278, 1.276, 1.275, 1.273, 1.271, 
    1.27, 1.269, 1.267, 1.266, 1.264, 1.263, 1.261, 1.26, 1.258, 1.257, 
    1.256, 1.254, 1.253, 1.251, 1.25, 1.248, 1.246, 1.245, 1.243, 1.241, 
    1.24, 1.238, 1.236, 1.234, 1.232, 1.231, 1.229, 1.227, 1.225, 1.223, 
    1.221, 1.219, 1.217, 1.214, 1.212, 1.21, 1.208, 1.205, 1.203, 1.201, 
    1.198, 1.195, 1.193, 1.19, 1.187, 1.185, 1.182, 1.179, 1.176, 1.173, 
    1.169, 1.166, 1.163, 1.159, 1.156, 1.152, 1.148, 1.145, 1.141, 1.137, 
    1.132, 1.128, 1.124, 1.119, 1.114, 1.109, 1.104, 1.099, 1.094, 1.088, 
    1.082, 1.076, 1.07, 1.063, 1.056, 1.049, 1.042, 1.034, 1.026, 1.018, 
    1.009, 1, 0.99, 0.98, 0.969, 0.957, 0.945, 0.933, 0.919, 0.905, 0.89, 
    0.874, 0.856, 0.838, 0.818, 0.797, 0.774, 0.75, 0.725, 0.699, 0.672, 
    0.645, 0.621, 0.6, 0.585, 0.577, 0.575, 0.579, 0.587, 0.601, 0.625, 
    0.663, 0.716, 0.777, 0.826, 0.844, 0.824, 0.779, 0.724, 0.671, 0.63, 
    0.605, 0.598, 0.609, 0.637, 0.684, 0.754, 0.851, 0.982, 1.153, 1.365, 
    1.601, 1.823, 1.986, 2.078, 2.126, 2.177, 2.259, 2.365, 2.458, 2.504, 
    2.501, 2.464, 2.409, 2.349, 2.289, 2.232, 2.179, 2.129, 2.084, 2.042, 
    2.003, 1.966, 1.932, 1.899, 1.868, 1.838, 1.809, 1.78, 1.752, 1.726, 
    1.706, 1.698, 1.713, 1.748, 1.777, 1.782, 1.769, 1.749, 1.727, 1.707, 
    1.692, 1.688, 1.695, 1.704, 1.705, 1.697, 1.682, 1.665, 1.648, 1.637, 
    1.642, 1.648, 1.639, 1.624, 1.61, 1.596, 1.583, 1.57, 1.558, 1.546, 
    1.533, 1.521, 1.51, 1.503, 1.505, 1.517, 1.527, 1.526, 1.518, 1.507, 
    1.495, 1.484, 1.474, 1.463, 1.453, 1.443, 1.433, 1.423, 1.412, 1.402, 
    1.392, 1.381, 1.37, 1.359, 1.347, 1.335, 1.323, 1.313, 1.308, 1.304, 
    1.294, 1.281, 1.266, 1.251, 1.235, 1.219, 1.203, 1.186, 1.169, 1.151, 
    1.133, 1.115, 1.097, 1.079, 1.062, 1.046, 1.031, 1.019, 1.009, 1.003, 
    0.999, 0.999, 1.001, 1.004, 1.007, 1.009, 1.008, 1.004, 0.999, 0.993, 
    0.992, 0.998, 1.018, 1.055, 1.109, 1.175, 1.247, 1.314, 1.383, 1.486, 
    1.674, 1.942, 2.143, 2.168, 2.08, 1.954, 1.817, 1.678, 1.538, 1.407, 
    1.315, 1.314, 1.451, 1.721, 2.019, 2.328, 2.744, 3.046, 3.073, 2.968, 
    2.843, 2.73, 2.634, 2.554, 2.486, 2.428, 2.379, 2.335, 2.297, 2.263, 
    2.233, 2.206, 2.181, 2.158 ;

 idx_rfr_montmorillonite_img = 0.001905461, 0.001659587, 0.002089296, 
    0.002187761, 0.002238721, 0.002570396, 0.002041738, 0.001949844, 
    0.001905461, 0.001174897, 0.0008317639, 0.0005888437, 0.0004677352, 
    0.0003548134, 0.0002511887, 0.0002041738, 0.0001230269, 0.0001071519, 
    5.248072e-05, 4.265796e-05, 3.388443e-05, 3.63078e-05, 4.466837e-05, 
    9.332538e-05, 9.772367e-05, 0.0001288249, 0.0001258925, 0.0001584893, 
    0.0001348963, 0.0001548817, 0.0001659587, 0.0001318256, 0.000245471, 
    0.0002344228, 0.0002187761, 0.0002630269, 0.0004073802, 0.0004570883, 
    0.0004365159, 0.000616595, 0.0007943284, 0.0007943284, 0.001380385, 
// NB: Relabel EgH79 value at 2.5 um as 2.4999 um to make room for 2.5 um Roush datum
// NB: Excise EgH79 value at 2.6 um in favor of Roush data
// end EgH79 Montmorillonite. Begin Roush Montmorillonite:
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.005, 0.005, 0.005, 0.006, 
    0.007, 0.008, 0.01, 0.013, 0.019, 0.028, 0.033, 0.025, 0.017, 0.012, 
    0.009, 0.008, 0.007, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 
    0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 
    0.006, 0.006, 0.006, 0.006, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 
    0.007, 0.007, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.01, 0.01, 0.01, 0.01, 0.01, 0.011, 0.011, 
    0.011, 0.011, 0.012, 0.012, 0.012, 0.013, 0.013, 0.013, 0.014, 0.014, 
    0.014, 0.015, 0.015, 0.015, 0.016, 0.016, 0.017, 0.017, 0.018, 0.018, 
    0.019, 0.02, 0.02, 0.021, 0.022, 0.023, 0.023, 0.024, 0.025, 0.026, 
    0.027, 0.028, 0.029, 0.031, 0.032, 0.034, 0.035, 0.037, 0.039, 0.041, 
    0.043, 0.045, 0.048, 0.05, 0.053, 0.057, 0.061, 0.065, 0.07, 0.075, 
    0.081, 0.088, 0.096, 0.105, 0.116, 0.129, 0.144, 0.163, 0.185, 0.212, 
    0.244, 0.282, 0.326, 0.375, 0.426, 0.478, 0.53, 0.582, 0.636, 0.691, 
    0.742, 0.78, 0.793, 0.774, 0.737, 0.706, 0.697, 0.718, 0.768, 0.841, 
    0.931, 1.03, 1.14, 1.25, 1.37, 1.49, 1.62, 1.74, 1.84, 1.9, 1.89, 1.82, 
    1.68, 1.54, 1.43, 1.37, 1.31, 1.22, 1.08, 0.919, 0.759, 0.623, 0.514, 
    0.43, 0.364, 0.313, 0.272, 0.24, 0.214, 0.193, 0.176, 0.162, 0.151, 
    0.142, 0.136, 0.132, 0.13, 0.133, 0.139, 0.152, 0.174, 0.204, 0.234, 
    0.242, 0.218, 0.183, 0.155, 0.136, 0.128, 0.128, 0.135, 0.145, 0.15, 
    0.141, 0.123, 0.106, 0.093, 0.086, 0.086, 0.093, 0.099, 0.086, 0.07, 
    0.06, 0.054, 0.051, 0.05, 0.049, 0.05, 0.051, 0.054, 0.059, 0.067, 0.078, 
    0.092, 0.097, 0.089, 0.075, 0.064, 0.057, 0.052, 0.05, 0.048, 0.047, 
    0.047, 0.047, 0.048, 0.049, 0.05, 0.051, 0.053, 0.055, 0.057, 0.06, 
    0.064, 0.068, 0.075, 0.083, 0.092, 0.093, 0.091, 0.092, 0.095, 0.1, 
    0.106, 0.113, 0.122, 0.131, 0.142, 0.155, 0.169, 0.186, 0.204, 0.225, 
    0.248, 0.274, 0.303, 0.334, 0.367, 0.401, 0.436, 0.47, 0.503, 0.535, 
    0.564, 0.594, 0.624, 0.657, 0.696, 0.743, 0.8, 0.866, 0.94, 1.02, 1.09, 
    1.15, 1.2, 1.24, 1.3, 1.38, 1.45, 1.4, 1.18, 0.921, 0.731, 0.621, 0.572, 
    0.572, 0.624, 0.739, 0.932, 1.19, 1.47, 1.66, 1.72, 1.75, 1.64, 1.27, 
    0.864, 0.592, 0.425, 0.321, 0.253, 0.206, 0.172, 0.147, 0.127, 0.112, 
    0.099, 0.089, 0.081, 0.073, 0.067, 0.062 ;
}

netcdf kaolinite_ior {
dimensions:
	bnd = 401 ;
variables:
	double bnd(bnd) ;
		bnd:units = "microns" ;
		bnd:longname = "band center wavelength" ;
		bnd:C_format = "%.5g" ;
	float idx_rfr_kaolinite_rl(bnd) ;
		idx_rfr_kaolinite_rl:units = "" ;
		idx_rfr_kaolinite_rl:longname = "kaolinite refractive index, real part " ;
		idx_rfr_kaolinite_rl:C_format = "%.4g" ;
	float idx_rfr_kaolinite_img(bnd) ;
		idx_rfr_kaolinite_img:units = "" ;
		idx_rfr_kaolinite_img:longname = "kaolinite refractive index, imag part " ;
		idx_rfr_kaolinite_img:C_format = "%.3g" ;

// global attributes:
		:description = "kaolinite refractive indices - T. Roush, Pollack, Orenberg, Icarus 94, 1991" ;
		:RCS_Header = "$Header: /home/zender/cvs/idx_rfr/roush/kaolinite_ior.cdl,v 1.1 2006-01-29 07:55:51 zender Exp $" ;
		:history = "" ;
		:author = "T. Roush(NASA Ames), Pollack, and Orenberg" ;
		:date = "netCDF file created 01 October, 2005" ;
data:

 bnd = 5, 5.01, 5.02, 5.03, 5.04, 5.05, 5.061, 5.071, 5.081, 5.092, 5.102, 
    5.113, 5.123, 5.134, 5.144, 5.155, 5.165, 5.176, 5.187, 5.198, 5.208, 
    5.219, 5.23, 5.241, 5.252, 5.263, 5.274, 5.285, 5.297, 5.308, 5.319, 
    5.331, 5.342, 5.353, 5.365, 5.376, 5.388, 5.4, 5.411, 5.423, 5.435, 
    5.447, 5.458, 5.47, 5.483, 5.495, 5.507, 5.519, 5.531, 5.543, 5.556, 
    5.568, 5.58, 5.593, 5.605, 5.618, 5.631, 5.643, 5.656, 5.669, 5.682, 
    5.695, 5.708, 5.721, 5.734, 5.747, 5.76, 5.774, 5.787, 5.8, 5.814, 5.827, 
    5.841, 5.855, 5.869, 5.882, 5.896, 5.91, 5.924, 5.938, 5.952, 5.967, 
    5.981, 5.995, 6.01, 6.024, 6.039, 6.053, 6.068, 6.083, 6.098, 6.113, 
    6.128, 6.142, 6.158, 6.173, 6.188, 6.203, 6.219, 6.234, 6.25, 6.266, 
    6.281, 6.297, 6.313, 6.329, 6.345, 6.361, 6.378, 6.394, 6.41, 6.427, 
    6.443, 6.46, 6.477, 6.494, 6.51, 6.527, 6.544, 6.562, 6.579, 6.596, 
    6.614, 6.631, 6.649, 6.667, 6.685, 6.702, 6.72, 6.739, 6.757, 6.775, 
    6.793, 6.812, 6.831, 6.849, 6.868, 6.887, 6.906, 6.925, 6.944, 6.964, 
    6.983, 7.003, 7.023, 7.042, 7.062, 7.082, 7.102, 7.122, 7.143, 7.163, 
    7.184, 7.205, 7.225, 7.246, 7.267, 7.289, 7.31, 7.331, 7.353, 7.375, 
    7.396, 7.418, 7.44, 7.463, 7.485, 7.508, 7.53, 7.553, 7.576, 7.599, 
    7.622, 7.645, 7.669, 7.692, 7.716, 7.74, 7.764, 7.788, 7.813, 7.837, 
    7.862, 7.886, 7.911, 7.937, 7.962, 7.987, 8.013, 8.039, 8.064, 8.091, 
    8.117, 8.143, 8.17, 8.197, 8.224, 8.251, 8.278, 8.306, 8.333, 8.361, 
    8.389, 8.417, 8.446, 8.475, 8.503, 8.532, 8.562, 8.591, 8.621, 8.651, 
    8.681, 8.711, 8.741, 8.772, 8.803, 8.834, 8.865, 8.897, 8.929, 8.961, 
    8.993, 9.025, 9.058, 9.091, 9.124, 9.158, 9.191, 9.225, 9.259, 9.294, 
    9.328, 9.363, 9.399, 9.434, 9.47, 9.506, 9.542, 9.578, 9.615, 9.653, 
    9.69, 9.728, 9.766, 9.804, 9.842, 9.881, 9.921, 9.96, 10, 10.04, 10.081, 
    10.121, 10.163, 10.204, 10.246, 10.288, 10.331, 10.373, 10.417, 10.46, 
    10.504, 10.549, 10.593, 10.638, 10.684, 10.73, 10.776, 10.823, 10.87, 
    10.917, 10.965, 11.013, 11.062, 11.111, 11.161, 11.211, 11.261, 11.312, 
    11.364, 11.416, 11.468, 11.521, 11.574, 11.628, 11.682, 11.737, 11.792, 
    11.848, 11.905, 11.962, 12.019, 12.077, 12.136, 12.195, 12.255, 12.315, 
    12.376, 12.438, 12.5, 12.563, 12.626, 12.69, 12.755, 12.821, 12.887, 
    12.953, 13.021, 13.089, 13.158, 13.228, 13.298, 13.369, 13.441, 13.514, 
    13.587, 13.661, 13.736, 13.812, 13.889, 13.966, 14.045, 14.124, 14.205, 
    14.286, 14.368, 14.451, 14.535, 14.62, 14.706, 14.793, 14.881, 14.97, 
    15.06, 15.152, 15.244, 15.337, 15.432, 15.528, 15.625, 15.723, 15.823, 
    15.924, 16.026, 16.129, 16.234, 16.34, 16.447, 16.556, 16.667, 16.779, 
    16.892, 17.007, 17.123, 17.241, 17.361, 17.483, 17.606, 17.731, 17.857, 
    17.986, 18.116, 18.248, 18.382, 18.519, 18.657, 18.797, 18.939, 19.084, 
    19.231, 19.38, 19.531, 19.685, 19.841, 20, 20.161, 20.325, 20.492, 
    20.661, 20.833, 21.008, 21.186, 21.368, 21.552, 21.739, 21.93, 22.124, 
    22.321, 22.523, 22.727, 22.936, 23.148, 23.364, 23.585, 23.81, 24.038, 
    24.272, 24.51, 24.752, 25 ;

 idx_rfr_kaolinite_rl = 1.362, 1.362, 1.362, 1.361, 1.361, 1.36, 1.36, 1.36, 
    1.359, 1.359, 1.358, 1.358, 1.357, 1.357, 1.357, 1.356, 1.356, 1.355, 
    1.355, 1.354, 1.354, 1.353, 1.353, 1.352, 1.352, 1.351, 1.351, 1.35, 
    1.35, 1.349, 1.349, 1.348, 1.348, 1.347, 1.347, 1.346, 1.346, 1.345, 
    1.345, 1.344, 1.343, 1.343, 1.342, 1.342, 1.341, 1.34, 1.34, 1.339, 
    1.339, 1.338, 1.337, 1.337, 1.336, 1.336, 1.335, 1.334, 1.334, 1.333, 
    1.332, 1.332, 1.331, 1.33, 1.329, 1.329, 1.328, 1.327, 1.327, 1.326, 
    1.325, 1.324, 1.324, 1.323, 1.322, 1.321, 1.32, 1.319, 1.319, 1.318, 
    1.317, 1.316, 1.315, 1.314, 1.314, 1.313, 1.312, 1.311, 1.31, 1.309, 
    1.308, 1.307, 1.306, 1.305, 1.304, 1.303, 1.302, 1.301, 1.3, 1.299, 
    1.298, 1.297, 1.296, 1.294, 1.293, 1.292, 1.291, 1.29, 1.288, 1.287, 
    1.286, 1.285, 1.283, 1.282, 1.281, 1.279, 1.278, 1.277, 1.275, 1.274, 
    1.272, 1.271, 1.269, 1.268, 1.266, 1.265, 1.263, 1.262, 1.26, 1.258, 
    1.256, 1.255, 1.253, 1.251, 1.249, 1.247, 1.245, 1.244, 1.242, 1.24, 
    1.237, 1.235, 1.233, 1.231, 1.229, 1.227, 1.224, 1.222, 1.22, 1.217, 
    1.215, 1.212, 1.21, 1.207, 1.204, 1.201, 1.199, 1.196, 1.193, 1.19, 
    1.187, 1.183, 1.18, 1.177, 1.173, 1.17, 1.166, 1.163, 1.159, 1.155, 
    1.151, 1.147, 1.142, 1.138, 1.133, 1.129, 1.124, 1.119, 1.114, 1.109, 
    1.103, 1.098, 1.092, 1.086, 1.08, 1.073, 1.066, 1.059, 1.052, 1.045, 
    1.037, 1.029, 1.02, 1.011, 1.002, 0.992, 0.981, 0.971, 0.959, 0.947, 
    0.934, 0.921, 0.906, 0.891, 0.874, 0.857, 0.837, 0.817, 0.794, 0.77, 
    0.743, 0.713, 0.68, 0.643, 0.601, 0.555, 0.506, 0.461, 0.433, 0.436, 
    0.479, 0.567, 0.669, 0.718, 0.685, 0.606, 0.514, 0.431, 0.37, 0.332, 
    0.312, 0.305, 0.308, 0.32, 0.34, 0.37, 0.411, 0.469, 0.549, 0.662, 0.825, 
    1.062, 1.397, 1.813, 2.184, 2.35, 2.304, 2.158, 2.065, 2.252, 2.692, 
    2.84, 2.714, 2.544, 2.393, 2.266, 2.157, 2.062, 1.975, 1.894, 1.817, 
    1.74, 1.661, 1.58, 1.503, 1.454, 1.494, 1.617, 1.676, 1.637, 1.615, 
    1.701, 1.803, 1.954, 2.217, 2.289, 2.218, 2.131, 2.056, 1.994, 1.942, 
    1.898, 1.86, 1.827, 1.796, 1.769, 1.744, 1.72, 1.698, 1.677, 1.657, 
    1.637, 1.619, 1.6, 1.582, 1.563, 1.545, 1.526, 1.506, 1.486, 1.465, 
    1.446, 1.435, 1.447, 1.481, 1.497, 1.487, 1.467, 1.443, 1.419, 1.396, 
    1.373, 1.355, 1.347, 1.359, 1.377, 1.377, 1.361, 1.339, 1.314, 1.289, 
    1.264, 1.239, 1.213, 1.187, 1.161, 1.136, 1.113, 1.093, 1.08, 1.076, 
    1.081, 1.092, 1.103, 1.105, 1.094, 1.07, 1.037, 1.003, 0.979, 0.98, 
    0.995, 0.983, 0.938, 0.882, 0.828, 0.784, 0.755, 0.742, 0.745, 0.76, 
    0.786, 0.818, 0.851, 0.881, 0.904, 0.924, 0.948, 0.987, 1.054, 1.159, 
    1.304, 1.476, 1.643, 1.783, 1.938, 2.234, 2.715, 3.071, 3.087, 2.936, 
    2.757, 2.59, 2.439, 2.3, 2.168, 2.039, 1.908, 1.77, 1.626, 1.493, 1.423, 
    1.505, 1.82, 2.368, 2.853, 2.973, 2.868, 2.709, 2.551, 2.405, 2.28, 2.21, 
    2.279, 2.535, 2.798, 2.879, 2.839, 2.765, 2.691, 2.625, 2.569, 2.52 ;

 idx_rfr_kaolinite_img = 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 0.005, 
    0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 0.005, 
    0.005, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 
    0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.008, 0.008, 0.008, 0.008, 
    0.008, 0.008, 0.009, 0.009, 0.009, 0.009, 0.01, 0.01, 0.01, 0.01, 0.011, 
    0.011, 0.011, 0.012, 0.012, 0.012, 0.013, 0.013, 0.013, 0.014, 0.014, 
    0.015, 0.015, 0.016, 0.016, 0.017, 0.018, 0.018, 0.019, 0.02, 0.021, 
    0.021, 0.022, 0.023, 0.024, 0.026, 0.027, 0.028, 0.03, 0.031, 0.033, 
    0.035, 0.038, 0.04, 0.043, 0.046, 0.05, 0.054, 0.059, 0.064, 0.071, 
    0.079, 0.089, 0.102, 0.119, 0.142, 0.174, 0.22, 0.287, 0.374, 0.475, 
    0.572, 0.636, 0.628, 0.553, 0.478, 0.448, 0.466, 0.525, 0.611, 0.708, 
    0.809, 0.911, 1.01, 1.12, 1.23, 1.35, 1.48, 1.62, 1.76, 1.93, 2.1, 2.26, 
    2.37, 2.34, 2.1, 1.74, 1.44, 1.31, 1.4, 1.58, 1.44, 0.979, 0.64, 0.454, 
    0.348, 0.284, 0.243, 0.215, 0.198, 0.189, 0.188, 0.195, 0.215, 0.254, 
    0.325, 0.443, 0.585, 0.638, 0.586, 0.574, 0.662, 0.761, 0.794, 0.856, 
    0.748, 0.483, 0.305, 0.21, 0.157, 0.124, 0.103, 0.089, 0.078, 0.071, 
    0.065, 0.06, 0.056, 0.053, 0.051, 0.05, 0.048, 0.048, 0.047, 0.047, 
    0.048, 0.049, 0.051, 0.054, 0.058, 0.065, 0.076, 0.095, 0.124, 0.156, 
    0.16, 0.134, 0.107, 0.091, 0.084, 0.083, 0.087, 0.098, 0.116, 0.14, 
    0.159, 0.154, 0.133, 0.116, 0.106, 0.102, 0.103, 0.107, 0.113, 0.122, 
    0.135, 0.151, 0.171, 0.195, 0.225, 0.258, 0.293, 0.323, 0.343, 0.35, 
    0.347, 0.341, 0.34, 0.35, 0.375, 0.417, 0.459, 0.472, 0.46, 0.46, 0.486, 
    0.535, 0.603, 0.682, 0.768, 0.855, 0.939, 1.02, 1.09, 1.15, 1.21, 1.27, 
    1.34, 1.43, 1.53, 1.66, 1.78, 1.88, 1.95, 1.98, 2, 2.08, 2.18, 2.09, 
    1.64, 1.16, 0.834, 0.637, 0.519, 0.446, 0.403, 0.383, 0.384, 0.407, 
    0.462, 0.564, 0.743, 1.02, 1.38, 1.72, 1.82, 1.5, 1.05, 0.732, 0.561, 
    0.485, 0.478, 0.541, 0.685, 0.885, 0.986, 0.844, 0.601, 0.415, 0.298, 
    0.224, 0.177, 0.144, 0.121 ;
}

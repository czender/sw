// ncgen -b -o ${DATA}/aca/idx_rfr_HKS98.nc ${HOME}/idx_rfr/idx_rfr_HKS98.cdl
// ncks -C -v idx_rfr_lac_HKS98_img,idx_rfr_lac_HKS98_rl ${DATA}/aca/idx_rfr_HKS98.nc
// scp ${DATA}/aca/idx_rfr_HKS98.nc dust.ess.uci.edu:/data/zender/aca

netcdf idx_rfr_HKS98 {
dimensions:
	bnd=62; // (62 currently)
variables:

// global attributes:

	:RCS_Header = "$Id$";
	:history = "";
	:description = "OPAC refractive indices" ;
	:source="
M. Hess and P. Koepke and I. Schult (1998) aka HKS98,
Optical Properties of Aerosols and Clouds: The Software Package OPAC,
Bull. Am. Meteorol. Soc, 79(5), 831--844

Homepage: http://www.lrz-muenchen.de/~uh234an/www/radaer/opac.html,
Software: ftp://ftp.lrz-muenchen.de/pub/science/meteorology/aerosol/opac/opac31a.tar.gz

File originally created with tbl2cdf from OPAC's soot00 file and waso?? files.

Note that most OPAC aerosol properties come from DKS91:
Atmospheric Aerosols: Global Climatology and Radiative Characteristics
by Guillaume A. d'Almeida and Peter Koepke and Eric P. Shettle

CSZ added channel at 0.2 microns to facilitate computation of dust optical properties in CCM spectral bands.
These data were copied from the HKS98 data at 0.25 microns if no other information was available.
There are now 62 bands.

20060601: MF added water soluble organic carbon (wsoc) refractive indecies from OPAC
          The two digits following 'wsoc' in the variable name are percent relative humidity.
20060604: CSZ changed soot to lac.";

	float bnd(bnd);
	bnd:long_name = "Band center wavelength";
	bnd:units = "micron";
	bnd:C_format = "%.5g";

	float idx_rfr_lac_HKS98_rl(bnd);
	idx_rfr_lac_HKS98_rl:long_name = "Light-absorbing carbon (soot) real index of refraction";
	idx_rfr_lac_HKS98_rl:units = "";
	idx_rfr_lac_HKS98_rl:C_format = "%.4g";

	float idx_rfr_lac_HKS98_img(bnd);
	idx_rfr_lac_HKS98_img:long_name = "Light-absorbing carbon (soot) imaginary index of refraction";
	idx_rfr_lac_HKS98_img:units = "";
	idx_rfr_lac_HKS98_img:C_format = "%.3g";

	float idx_rfr_wsoc00_HKS98_rl(bnd);
	idx_rfr_wsoc00_HKS98_rl:long_name = "Water soluble organic/inorganic mixture real index of refraction";
	idx_rfr_wsoc00_HKS98_rl:units = "";
	idx_rfr_wsoc00_HKS98_rl:C_format = "%.4g";

	float idx_rfr_wsoc00_HKS98_img(bnd);
	idx_rfr_wsoc00_HKS98_img:long_name = "Water soluble organic/inorganic mixture imaginary index of refraction, dry";
	idx_rfr_wsoc00_HKS98_img:units = "";
	idx_rfr_wsoc00_HKS98_img:C_format = "%.3g";

	float idx_rfr_wsoc50_HKS98_rl(bnd);
	idx_rfr_wsoc50_HKS98_rl:long_name = "Water soluble organic/inorganic mixture real index of refraction, RH=0.50";
	idx_rfr_wsoc50_HKS98_rl:units = "";
	idx_rfr_wsoc50_HKS98_rl:C_format = "%.4g";

	float idx_rfr_wsoc50_HKS98_img(bnd);
	idx_rfr_wsoc50_HKS98_img:long_name = "Water soluble organic/inorganic mixture imaginary index of refraction, RH=0.50";
	idx_rfr_wsoc50_HKS98_img:units = "";
	idx_rfr_wsoc50_HKS98_img:C_format = "%.3g";

	float idx_rfr_wsoc70_HKS98_rl(bnd);
	idx_rfr_wsoc70_HKS98_rl:long_name = "Water soluble organic/inorganic mixture real index of refraction, RH=0.70";
	idx_rfr_wsoc70_HKS98_rl:units = "";
	idx_rfr_wsoc70_HKS98_rl:C_format = "%.4g";

	float idx_rfr_wsoc70_HKS98_img(bnd);
	idx_rfr_wsoc70_HKS98_img:long_name = "Water soluble organic/inorganic mixture imaginary index of refraction, RH=0.70";
	idx_rfr_wsoc70_HKS98_img:units = "";
	idx_rfr_wsoc70_HKS98_img:C_format = "%.3g";

	float idx_rfr_wsoc80_HKS98_rl(bnd);
	idx_rfr_wsoc80_HKS98_rl:long_name = "Water soluble organic/inorganic mixture real index of refraction, RH=0.80";
	idx_rfr_wsoc80_HKS98_rl:units = "";
	idx_rfr_wsoc80_HKS98_rl:C_format = "%.4g";

	float idx_rfr_wsoc80_HKS98_img(bnd);
	idx_rfr_wsoc80_HKS98_img:long_name = "Water soluble organic/inorganic mixture imaginary index of refraction, RH=0.80";
	idx_rfr_wsoc80_HKS98_img:units = "";
	idx_rfr_wsoc80_HKS98_img:C_format = "%.3g";

	float idx_rfr_wsoc90_HKS98_rl(bnd);
	idx_rfr_wsoc90_HKS98_rl:long_name = "Water soluble organic/inorganic mixture real index of refraction, RH=0.90";
	idx_rfr_wsoc90_HKS98_rl:units = "";
	idx_rfr_wsoc90_HKS98_rl:C_format = "%.4g";

	float idx_rfr_wsoc90_HKS98_img(bnd);
	idx_rfr_wsoc90_HKS98_img:long_name = "Water soluble organic/inorganic mixture imaginary index of refraction, RH=0.90";
	idx_rfr_wsoc90_HKS98_img:units = "";
	idx_rfr_wsoc90_HKS98_img:C_format = "%.3g";

	float idx_rfr_wsoc95_HKS98_rl(bnd);
	idx_rfr_wsoc95_HKS98_rl:long_name = "Water soluble organic/inorganic mixture real index of refraction, RH=0.95";
	idx_rfr_wsoc95_HKS98_rl:units = "";
	idx_rfr_wsoc95_HKS98_rl:C_format = "%.4g";

	float idx_rfr_wsoc95_HKS98_img(bnd);
	idx_rfr_wsoc95_HKS98_img:long_name = "Water soluble organic/inorganic mixture imaginary index of refraction, RH=0.95";
	idx_rfr_wsoc95_HKS98_img:units = "";
	idx_rfr_wsoc95_HKS98_img:C_format = "%.3g";

	float idx_rfr_wsoc98_HKS98_rl(bnd);
	idx_rfr_wsoc98_HKS98_rl:long_name = "Water soluble organic/inorganic mixture real index of refraction, RH=0.98";
	idx_rfr_wsoc98_HKS98_rl:units = "";
	idx_rfr_wsoc98_HKS98_rl:C_format = "%.4g";

	float idx_rfr_wsoc98_HKS98_img(bnd);
	idx_rfr_wsoc98_HKS98_img:long_name = "Water soluble organic/inorganic mixture imaginary index of refraction, RH=0.98";
	idx_rfr_wsoc98_HKS98_img:units = "";
	idx_rfr_wsoc98_HKS98_img:C_format = "%.3g";

	float idx_rfr_wsoc99_HKS98_rl(bnd);
	idx_rfr_wsoc99_HKS98_rl:long_name = "Water soluble organic/inorganic mixture real index of refraction, RH=0.99";
	idx_rfr_wsoc99_HKS98_rl:units = "";
	idx_rfr_wsoc99_HKS98_rl:C_format = "%.4g";

	float idx_rfr_wsoc99_HKS98_img(bnd);
	idx_rfr_wsoc99_HKS98_img:long_name = "Water soluble organic/inorganic mixture imaginary index of refraction, RH=0.99";
	idx_rfr_wsoc99_HKS98_img:units = "";
	idx_rfr_wsoc99_HKS98_img:C_format = "%.3g";

data:

 bnd = 0.20, 0.25, 0.3, 0.35, 0.4, 0.45, 0.5, 0.55, 0.6, 0.65, 0.7, 0.75, 0.8, 0.9, 
    1, 1.25, 1.5, 1.75, 2, 2.5, 3, 3.2, 3.39, 3.5, 3.75, 4, 4.5, 5, 5.5, 6, 
    6.2, 6.5, 7.2, 7.9, 8.2, 8.5, 8.7, 9, 9.2, 9.5, 9.8, 10, 10.6, 11, 11.5, 
    12.5, 13, 14, 14.8, 15, 16.4, 17.2, 18, 18.5, 20, 21.3, 22.5, 25, 27.9, 
    30, 35, 40 ;

 idx_rfr_lac_HKS98_rl = 1.62, 1.62, 1.74, 1.75, 1.75, 1.75, 1.75, 1.75, 1.75, 
    1.75, 1.75, 1.75, 1.75, 1.75, 1.76, 1.76, 1.77, 1.79, 1.8, 1.82, 1.84, 
    1.86, 1.87, 1.88, 1.9, 1.92, 1.94, 1.97, 1.99, 2.02, 2.03, 2.04, 2.06, 
    2.12, 2.13, 2.15, 2.16, 2.17, 2.18, 2.19, 2.2, 2.21, 2.22, 2.23, 2.24, 
    2.27, 2.28, 2.31, 2.33, 2.33, 2.36, 2.38, 2.4, 2.41, 2.45, 2.46, 2.48, 
    2.51, 2.54, 2.57, 2.63, 2.69 ;

 idx_rfr_lac_HKS98_img = 0.45, 0.45, 0.47, 0.465, 0.46, 0.455, 0.45, 0.44, 
    0.435, 0.435, 0.43, 0.43, 0.43, 0.435, 0.44, 0.45, 0.46, 0.48, 
    0.49, 0.51, 0.54, 0.54, 0.5495, 0.56, 0.57, 0.58, 0.59, 0.6, 
    0.61, 0.62, 0.625, 0.63, 0.65, 0.67, 0.68, 0.69, 0.69, 0.7, 
    0.7, 0.71, 0.715, 0.72, 0.73, 0.73, 0.74, 0.75, 0.76, 0.775, 
    0.79, 0.79, 0.81, 0.82, 0.825, 0.83, 0.85, 0.86, 0.87, 0.89, 
    0.91, 0.93, 0.97, 1 ;


 idx_rfr_wsoc00_HKS98_rl = 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53,
    1.52, 1.52, 1.52, 1.51, 1.51, 1.47, 1.42, 1.42, 1.42, 1.43, 1.43, 1.45,
    1.452, 1.455, 1.46, 1.45, 1.44, 1.41, 1.43, 1.46, 1.4, 1.2, 1.01, 1.3,
    2.4, 2.56, 2.2, 1.95, 1.87, 1.82, 1.76, 1.72, 1.67, 1.62, 1.62, 1.56,
    1.44, 1.42, 1.75, 2.08, 1.98, 1.85, 2.12, 2.06, 2, 1.88, 1.84, 1.82,
    1.92, 1.86 ;

 idx_rfr_wsoc00_HKS98_img = 0.03, 0.03, 0.008, 0.005, 0.005, 0.005, 0.005, 0.006, 0.006, 0.007,
    0.007, 0.0085, 0.01, 0.013, 0.0155, 0.019, 0.0225, 0.0175, 0.008, 0.012,
    0.022, 0.008, 0.00705, 0.005, 0.004, 0.005, 0.013, 0.012, 0.018, 0.023,
    0.027, 0.033, 0.07, 0.065, 0.1, 0.215, 0.29, 0.37, 0.42, 0.16, 0.095,
    0.09, 0.07, 0.05, 0.047, 0.053, 0.055, 0.073, 0.1, 0.2, 0.16, 0.242,
    0.18, 0.17, 0.22, 0.23, 0.24, 0.28, 0.29, 0.3, 0.4, 0.5 ;


 idx_rfr_wsoc50_HKS98_rl = 1.451, 1.451, 1.445, 1.442, 1.44, 1.439, 1.438, 1.437, 1.437, 1.436,
    1.436, 1.436, 1.43, 1.43, 1.429, 1.422, 1.421, 1.396, 1.366, 1.345,
    1.397, 1.453, 1.427, 1.426, 1.413, 1.406, 1.4, 1.391, 1.373, 1.342,
    1.398, 1.403, 1.359, 1.244, 1.14, 1.29, 1.87, 1.95, 1.756, 1.618, 1.569,
    1.537, 1.487, 1.453, 1.414, 1.386, 1.397, 1.395, 1.354, 1.349, 1.56,
    1.754, 1.718, 1.659, 1.819, 1.792, 1.768, 1.716, 1.703, 1.694, 1.738, 1.7 ;

 idx_rfr_wsoc50_HKS98_img = 0.01589, 0.01589, 0.004238, 0.002649, 0.002649, 0.002649, 0.002649,
    0.003179, 0.003179, 0.003709, 0.003709, 0.004503, 0.005298, 0.006887,
    0.008213, 0.01007, 0.01201, 0.009318, 0.004756, 0.007176, 0.1396,
    0.04769, 0.01462, 0.007069, 0.003765, 0.004812, 0.01319, 0.01219,
    0.01499, 0.0625, 0.05568, 0.03592, 0.05218, 0.05038, 0.06948, 0.1312,
    0.1715, 0.2148, 0.242, 0.1056, 0.07285, 0.07157, 0.06878, 0.07201,
    0.09167, 0.1499, 0.1726, 0.2127, 0.2392, 0.295, 0.2855, 0.3299, 0.2957,
    0.288, 0.3013, 0.3001, 0.3011, 0.3157, 0.313, 0.3132, 0.3699, 0.4459 ;


 idx_rfr_wsoc70_HKS98_rl = 1.431, 1.431, 1.423, 1.42, 1.418, 1.416, 1.415, 1.414, 1.413, 1.413,
    1.413, 1.412, 1.408, 1.407, 1.406, 1.4, 1.399, 1.378, 1.353, 1.326,
    1.391, 1.458, 1.426, 1.421, 1.403, 1.394, 1.385, 1.376, 1.356, 1.325,
    1.391, 1.389, 1.348, 1.255, 1.172, 1.287, 1.736, 1.796, 1.644, 1.534,
    1.493, 1.466, 1.418, 1.386, 1.35, 1.328, 1.341, 1.354, 1.333, 1.332,
    1.512, 1.672, 1.652, 1.611, 1.743, 1.725, 1.709, 1.675, 1.669, 1.662,
    1.692, 1.659 ;

 idx_rfr_wsoc70_HKS98_img = 0.01235, 0.01235, 0.003293, 0.002058, 0.002058, 0.002058, 0.002058,
    0.00247, 0.00247, 0.002881, 0.002881, 0.003499, 0.004116, 0.005351,
    0.006381, 0.007825, 0.009379, 0.007262, 0.00394, 0.005963, 0.1691,
    0.05766, 0.01652, 0.007589, 0.003706, 0.004765, 0.01324, 0.01224,
    0.01423, 0.07243, 0.06289, 0.03665, 0.0477, 0.0467, 0.06181, 0.1101,
    0.1417, 0.1758, 0.1973, 0.09198, 0.06729, 0.06693, 0.06847, 0.07754,
    0.1029, 0.1742, 0.2021, 0.2478, 0.2742, 0.3189, 0.3171, 0.352, 0.3247,
    0.3177, 0.3218, 0.3177, 0.3165, 0.3247, 0.3188, 0.3165, 0.3623, 0.4323 ;


 idx_rfr_wsoc80_HKS98_rl = 1.418, 1.418, 1.409, 1.405, 1.403, 1.401, 1.4, 1.399, 1.398, 1.397,
    1.397, 1.397, 1.393, 1.392, 1.391, 1.385, 1.384, 1.365, 1.344, 1.314,
    1.387, 1.462, 1.425, 1.417, 1.397, 1.386, 1.375, 1.367, 1.345, 1.313,
    1.385, 1.379, 1.341, 1.263, 1.194, 1.285, 1.647, 1.694, 1.569, 1.478,
    1.442, 1.418, 1.372, 1.342, 1.307, 1.288, 1.304, 1.326, 1.319, 1.32,
    1.48, 1.617, 1.608, 1.578, 1.693, 1.68, 1.67, 1.647, 1.646, 1.64, 1.661,
    1.632 ;

 idx_rfr_wsoc80_HKS98_img = 0.009976, 0.009976, 0.00266, 0.001663, 0.001663, 0.001663, 0.001663,
    0.001995, 0.001995, 0.002328, 0.002328, 0.002827, 0.003325, 0.004323,
    0.005156, 0.006324, 0.007616, 0.005886, 0.003395, 0.005152, 0.1889,
    0.06433, 0.01779, 0.007937, 0.003666, 0.004733, 0.01327, 0.01227,
    0.01373, 0.07907, 0.06772, 0.03714, 0.0447, 0.04424, 0.05668, 0.09599,
    0.1217, 0.1497, 0.1674, 0.08284, 0.06356, 0.06384, 0.06826, 0.08124,
    0.1104, 0.1905, 0.2219, 0.2712, 0.2976, 0.3348, 0.3382, 0.3668, 0.3442,
    0.3375, 0.3355, 0.3295, 0.3268, 0.3307, 0.3227, 0.3187, 0.3573, 0.4232 ;


 idx_rfr_wsoc90_HKS98_rl = 1.4, 1.4, 1.39, 1.385, 1.382, 1.381, 1.379, 1.378, 1.377, 1.376,
    1.376, 1.375, 1.372, 1.371, 1.371, 1.365, 1.364, 1.348, 1.332, 1.297,
    1.382, 1.467, 1.425, 1.411, 1.388, 1.375, 1.361, 1.353, 1.33, 1.298,
    1.378, 1.366, 1.332, 1.273, 1.224, 1.283, 1.527, 1.555, 1.469, 1.403,
    1.374, 1.354, 1.31, 1.281, 1.249, 1.235, 1.253, 1.289, 1.299, 1.304,
    1.437, 1.543, 1.549, 1.535, 1.625, 1.62, 1.618, 1.61, 1.615, 1.612, 1.62,
    1.596 ;

 idx_rfr_wsoc90_HKS98_img = 0.006783, 0.006783, 0.001809, 0.00113, 0.00113, 0.00113, 0.00113,
    0.001357, 0.001357, 0.001583, 0.001583, 0.001922, 0.002261, 0.002939,
    0.003507, 0.004302, 0.005242, 0.004034, 0.00266, 0.00406, 0.2155,
    0.07332, 0.01951, 0.008405, 0.003613, 0.00469, 0.01331, 0.01231, 0.01305,
    0.08801, 0.07421, 0.0378, 0.04067, 0.04093, 0.04977, 0.07701, 0.0949,
    0.1145, 0.1271, 0.07054, 0.05855, 0.05966, 0.06799, 0.08622, 0.1205,
    0.2124, 0.2485, 0.3029, 0.3291, 0.3563, 0.3666, 0.3867, 0.3704, 0.3643,
    0.3539, 0.3453, 0.3406, 0.3388, 0.3279, 0.3217, 0.3505, 0.411 ;


 idx_rfr_wsoc95_HKS98_rl = 1.387, 1.387, 1.376, 1.371, 1.368, 1.366, 1.364, 1.363, 1.362, 1.361,
    1.361, 1.36, 1.358, 1.357, 1.356, 1.351, 1.349, 1.337, 1.323, 1.285,
    1.378, 1.471, 1.424, 1.407, 1.381, 1.367, 1.351, 1.344, 1.319, 1.287,
    1.373, 1.357, 1.325, 1.28, 1.245, 1.281, 1.441, 1.457, 1.397, 1.349,
    1.325, 1.308, 1.266, 1.238, 1.208, 1.198, 1.217, 1.262, 1.285, 1.292,
    1.407, 1.49, 1.507, 1.504, 1.576, 1.576, 1.58, 1.583, 1.593, 1.591, 1.59,
    1.57 ;

 idx_rfr_wsoc95_HKS98_img = 0.0045, 0.0045, 0.0012, 0.00075, 0.00075, 0.00075, 0.00075, 0.0009,
    0.0009, 0.00105, 0.00105, 0.001275, 0.0015, 0.00195, 0.002327, 0.002857,
    0.003545, 0.00271, 0.002135, 0.003279, 0.2345, 0.07974, 0.02073, 0.00874,
    0.003575, 0.00466, 0.01334, 0.01234, 0.01256, 0.0944, 0.07885, 0.03827,
    0.03778, 0.03856, 0.04483, 0.06344, 0.07571, 0.08941, 0.09827, 0.06174,
    0.05496, 0.05668, 0.06779, 0.08978, 0.1278, 0.2281, 0.2675, 0.3255,
    0.3516, 0.3717, 0.387, 0.401, 0.3891, 0.3834, 0.3671, 0.3567, 0.3505,
    0.3446, 0.3317, 0.3238, 0.3456, 0.4022 ;


 idx_rfr_wsoc98_HKS98_rl = 1.377, 1.377, 1.365, 1.36, 1.356, 1.354, 1.352, 1.35, 1.349, 1.349,
    1.349, 1.348, 1.346, 1.345, 1.344, 1.34, 1.338, 1.327, 1.316, 1.275,
    1.375, 1.474, 1.424, 1.404, 1.376, 1.36, 1.343, 1.336, 1.311, 1.278,
    1.369, 1.35, 1.32, 1.286, 1.262, 1.28, 1.372, 1.377, 1.338, 1.305, 1.286,
    1.271, 1.23, 1.203, 1.174, 1.167, 1.188, 1.241, 1.274, 1.283, 1.382,
    1.447, 1.472, 1.479, 1.537, 1.541, 1.55, 1.562, 1.575, 1.575, 1.566, 1.549 ;

 idx_rfr_wsoc98_HKS98_img = 0.00265, 0.00265, 0.0007068, 0.0004417, 0.0004417, 0.0004417, 0.0004417,
    0.0005301, 0.0005301, 0.0006184, 0.0006185, 0.0007511, 0.0008836,
    0.001149, 0.001372, 0.001687, 0.00217, 0.001637, 0.00171, 0.002646,
    0.2499, 0.08494, 0.02172, 0.009011, 0.003544, 0.004635, 0.01336, 0.01236,
    0.01217, 0.09958, 0.08261, 0.03865, 0.03545, 0.03665, 0.04083, 0.05245,
    0.06017, 0.06906, 0.07494, 0.05461, 0.05206, 0.05426, 0.06763, 0.09267,
    0.1336, 0.2408, 0.2829, 0.3438, 0.3698, 0.3842, 0.4034, 0.4125, 0.4043,
    0.3988, 0.3777, 0.3658, 0.3585, 0.3493, 0.3347, 0.3255, 0.3417, 0.3952 ;


 idx_rfr_wsoc99_HKS98_rl = 1.373, 1.373, 1.36, 1.355, 1.351, 1.349, 1.347, 1.345, 1.344, 1.343,
    1.343, 1.343, 1.341, 1.34, 1.339, 1.335, 1.333, 1.323, 1.313, 1.271,
    1.374, 1.475, 1.423, 1.403, 1.374, 1.358, 1.34, 1.333, 1.307, 1.274,
    1.367, 1.347, 1.318, 1.288, 1.269, 1.279, 1.343, 1.343, 1.314, 1.287,
    1.269, 1.256, 1.215, 1.188, 1.16, 1.154, 1.176, 1.232, 1.269, 1.279,
    1.371, 1.429, 1.458, 1.468, 1.52, 1.527, 1.537, 1.553, 1.567, 1.568,
    1.556, 1.54 ;

 idx_rfr_wsoc99_HKS98_img = 0.001877, 0.001877, 0.0005006, 0.0003129, 0.0003129, 0.0003129, 0.0003129,
    0.0003754, 0.0003754, 0.000438, 0.000438, 0.000532, 0.0006258, 0.0008139,
    0.0009726, 0.001197, 0.001595, 0.001189, 0.001532, 0.002382, 0.2564,
    0.08712, 0.02214, 0.009125, 0.003531, 0.004625, 0.01337, 0.01237, 0.012,
    0.1017, 0.08418, 0.03881, 0.03447, 0.03585, 0.03916, 0.04786, 0.05367,
    0.06056, 0.06518, 0.05163, 0.05085, 0.05325, 0.06756, 0.09387, 0.1361,
    0.2461, 0.2894, 0.3514, 0.3775, 0.3894, 0.4103, 0.4173, 0.4106, 0.4053,
    0.3822, 0.3697, 0.3619, 0.3512, 0.3359, 0.3262, 0.34, 0.3922 ;

}

// ncgen -b -o $DATA/aca/idx_rfr_DKS91.nc $HOME/idx_rfr/idx_rfr_DKS91.cdl
// ncks -C -H -v idx_rfr_mineral_dust_img,idx_rfr_mineral_dust_rl $DATA/aca/idx_rfr_DKS91.nc

netcdf idx_rfr_DKS91 {
dimensions:
	bnd=62;
variables:

	:RCS_Header = "$Id$";
	:history = "";
	:source="Atmospheric Aerosols: Global Climatology and Radiative Characteristics
by Guillaume A. d'Almeida and Peter Koepke and Eric P. Shettle
Table 4.3, pp. 57-59, entered by CSZ 96/07/25

Mon Oct 13 11:25:43 MDT 1997: 
Added channels at 0.2 and 0.25 microns to facilitate computation of dust optical properties in CCM spectral bands.
These data were copied from the DKS91 data at 0.3 microns if no other information was available.
Indices from compilation of Shettle (from HITRAN96 CDROM) for Dust-like aerosol were used for 0.2 and 0.25 micron bands for both mineral_dust and dust_like aerosols.
NB: dust_like aerosol is MUCH weaker optically than Saharan dust in IR.
Indices from compilation of Shettle (from HITRAN96 CDROM) for H2SO4 at 300K (from HITRAN96 CDROM) were used for 0.2 and 0.25 micron bands for sulfate.
There are now 62 bands.";

	float bnd(bnd);
	bnd:long_name = "Band center wavelength";
	bnd:units = "micron";
	bnd:C_format = "%.5g";

	float idx_rfr_dust_like_rl(bnd);
	idx_rfr_dust_like_rl:long_name = "Dust-like real index of refraction";
	idx_rfr_dust_like_rl:units = "";
	idx_rfr_dust_like_rl:C_format = "%.4g";

	float idx_rfr_dust_like_img(bnd);
	idx_rfr_dust_like_img:long_name = "Dust-like imaginary index of refraction";
	idx_rfr_dust_like_img:units = "";
	idx_rfr_dust_like_img:C_format = "%.3g";

	float idx_rfr_mineral_dust_rl(bnd);
	idx_rfr_mineral_dust_rl:long_name = "Mineral dust real index of refraction";
	idx_rfr_mineral_dust_rl:units = "";
	idx_rfr_mineral_dust_rl:C_format = "%.4g";

	float idx_rfr_mineral_dust_img(bnd);
	idx_rfr_mineral_dust_img:long_name = "Mineral dust imaginary index of refraction";
	idx_rfr_mineral_dust_img:units = "";
	idx_rfr_mineral_dust_img:C_format = "%.3g";

	float idx_rfr_sulfate_rl(bnd);
	idx_rfr_sulfate_rl:long_name = "Sulfate real index of refraction";
	idx_rfr_sulfate_rl:units = "";
	idx_rfr_sulfate_rl:C_format = "%.4g";

	float idx_rfr_sulfate_img(bnd);
	idx_rfr_sulfate_img:long_name = "Sulfate imaginary index of refraction";
	idx_rfr_sulfate_img:units = "";
	idx_rfr_sulfate_img:C_format = "%.3g";

data:	
 bnd = 0.2, 0.25,
    0.3, 0.35, 0.4, 0.45, 0.5, 0.55, 0.6, 0.65, 0.7, 0.75, 0.8, 
    0.9, 1, 1.25, 1.5, 1.75, 2, 2.5, 3, 3.2, 3.392, 3.5, 3.75, 4, 4.5, 5, 
    5.5, 6, 6.2, 6.5, 7.2, 7.9, 8.2, 8.5, 8.7, 9, 9.2, 9.5, 9.8, 10, 10.951, 
    11, 11.5, 12.5, 13, 14, 14.8, 15, 16.4, 17.2, 18, 18.5, 20, 21.3, 22.5, 
    25, 27.9, 30, 35, 40 ;
 
 idx_rfr_dust_like_rl = 1.53, 1.53,
    1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 
    1.53, 1.52, 1.52, 1.52, 1.46, 1.41, 1.34, 1.26, 1.18, 1.16, 1.22, 1.26, 
    1.28, 1.27, 1.26, 1.26, 1.25, 1.22, 1.15, 1.14, 1.13, 1.4, 1.15, 1.13, 
    1.3, 1.4, 1.7, 1.72, 1.73, 1.74, 1.75, 1.62, 1.62, 1.59, 1.51, 1.47, 
    1.52, 1.57, 1.57, 1.6, 1.63, 1.64, 1.64, 1.68, 1.77, 1.9, 1.97, 1.89, 
    1.8, 1.9, 2.1 ;
 
 idx_rfr_dust_like_img = 0.070, 0.030,
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.009, 
    0.012, 0.01, 0.013, 0.011, 0.011, 0.012, 0.014, 0.016, 0.021, 0.037, 
    0.039, 0.042, 0.055, 0.04, 0.0742, 0.09, 0.1, 0.14, 0.15, 0.162, 0.162, 
    0.162, 0.12, 0.105, 0.1, 0.09, 0.1, 0.085, 0.01, 0.1, 0.1, 0.1, 0.115, 
    0.12, 0.22, 0.28, 0.28, 0.244, 0.32, 0.42, 0.5, 0.6 ;

 idx_rfr_mineral_dust_rl = 1.53, 1.53,
    1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 
    1.53, 1.53, 1.53, 1.53, 1.53, 1.42, 1.37, 1.267, 1.18, 1.16, 1.22, 1.26, 
    1.28, 1.27, 1.26, 1.26, 1.25, 1.22, 1.22, 1.14, 1.13, 1.4, 1.15, 1.13, 
    1.3, 1.4, 1.4, 1.72, 1.73, 1.74, 1.75, 1.30, 1.62, 1.59, 1.51, 1.47, 
    1.52, 1.57, 1.57, 1.6, 1.63, 1.64, 1.64, 1.68, 1.77, 1.9, 1.97, 1.89, 
    1.8, 1.9, 2.1 ;
 
 idx_rfr_mineral_dust_img = 0.070, 0.030, 
    2.5e-2, 1.70e-2, 1.30e-2, 8.50e-3, 7.80e-3, 5.50e-3, 4.50e-3, 4.50e-3, 
    4.00e-3, 4.00e-3, 1.20e-3, 1.20e-3, 1.00e-3, 1.30e-3, 1.40e-3, 1.80e-3, 2.00e-3, 3.40e-3, 
    0.012, 0.01, 0.013, 0.011, 0.011, 0.012, 0.014, 0.016, 0.021, 2.1e-2, 
    0.039, 0.042, 0.055, 0.04, 0.0742, 0.09, 0.1, 0.14, 0.15, 0.162, 0.162, 
    0.162, 9.e-2, 0.105, 0.1, 0.09, 0.1, 0.085, 0.01, 0.1, 0.1, 0.1, 0.115, 
    0.12, 0.22, 0.28, 0.28, 0.244, 0.32, 0.42, 0.5, 0.6 ;

 idx_rfr_sulfate_rl = 1.498, 1.484, 
    1.469, 1.452, 1.44, 1.432, 1.431, 1.43, 1.429, 1.429, 
    1.428, 1.427, 1.426, 1.425, 1.423, 1.41, 1.403, 1.39, 1.384, 1.344, 
    1.293, 1.311, 1.352, 1.376, 1.396, 1.398, 1.385, 1.36, 1.337, 1.425, 
    1.424, 1.37, 1.21, 1.14, 1.2, 1.37, 1.53, 1.65, 1.6, 1.67, 1.91, 1.89, 
    1.72, 1.67, 1.89, 1.74, 1.69, 1.64, 1.61, 1.59, 1.52, 1.724, 1.95, 1.927, 
    1.823, 1.78, 1.87, 1.93, 1.92, 1.92, 1.9, 1.89 ;
 
 idx_rfr_sulfate_img = 1e-08, 1e-08,
    1e-08, 1e-08, 1e-08, 1e-08, 1e-08, 1e-08, 1.47e-08, 
    1.47e-08, 1.99e-08, 1.89e-08, 1.7e-08, 1.79e-07, 1.5e-06, 1e-05, 
    0.000134, 0.00055, 0.00126, 0.00376, 0.0955, 0.135, 0.159, 0.158, 0.131, 
    0.136, 0.12, 0.121, 0.183, 0.195, 0.165, 0.128, 0.176, 0.488, 0.645, 
    0.755, 0.772, 0.633, 0.586, 0.75, 0.68, 0.455, 0.34, 0.485, 0.374, 0.198, 
    0.195, 0.195, 0.205, 0.211, 0.414, 0.59, 0.041, 0.0302, 0.0235, 0.292, 
    0.0315, 0.2, 0.18, 0.18, 0.19, 0.22 ;
}

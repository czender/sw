// $Id$
// ncgen -b -o ${DATA}/aca/idx_rfr_roush_illite.nc ${HOME}/idx_rfr/idx_rfr_roush_illite.cdl

netcdf idx_rfr_roush_illite {
dimensions:
	bnd = 3951 ;
	bnd_EgH79 = 44 ;

variables:

// global attributes:
	:RCS_Header = "$Id$" ;
	:history = "" ;
	:description = "Illite refractive indices" ;
	:source="
Ted Roush (NASA Ames) <troush at mail dot arc dot nasa dot gov>
Brian Hansell (UCLA) converted Roush's IR data into netCDF format 01 October, 2005.
Charlie Zender (UCI) <zender at uci dot edu> standardized 20060129.

Changed coordinate from wavenumber to wavelength.
Measured by Marvin Querry and reported in 1987 U.S. Army tech. note CRDEC-CR-88009
from Aberdeen, MD.

Begin Original e-mail header accompanying data from T. Roush:
From:	IO::memilham@CRDEC-VAX4.ARPA 14-JUN-1988 04:35
To:	HAL::DALTON
Subj:	Optical Constants: Illite

Received: from CRDEC-VAX4.ARPA by ames-io.ARPA with INTERNET ;
          Tue, 14 Jun 88 04:26:36 PDT
Date:     Tue, 14 Jun 88 7:23:56 EDT
From:     Merrill E. Milham <memilham@CRDEC-VAX4.ARPA>
To:       dalton%hal@AMES-IO.ARPA
Subject:  Optical Constants: Illite
Message-ID:  <8806140723.aa24544@CRDEC-VAX4.CRDEC-VAX4.ARPA>
Date:     Wed, 27 May 87 13:24 CDT
Subject:  OPT. CON. OF ILLITE WITH FIR DATA
To:       MEMILHAM@CRDEC.ARPA QUERRY
End Original e-mail header accompanying data from T. Roush
	";

	float bnd(bnd) ;
		bnd:units = "microns" ;
		bnd:longname = "Band center wavelength" ;
		bnd:C_format = "%.5g" ;

	float bnd_wvn(bnd) ;
		bnd_wvn:units = "cm-1" ;
		bnd_wvn:longname = "Band center wavenumber" ;
		bnd_wvn:C_format = "%.5g" ;

	float idx_rfr_illite_rl(bnd) ;
		idx_rfr_illite_rl:units = "" ;
		idx_rfr_illite_rl:longname = "Illite refractive index, real part " ;
		idx_rfr_illite_rl:C_format = "%.4g" ;

	float idx_rfr_illite_img(bnd) ;
		idx_rfr_illite_img:units = "" ;
		idx_rfr_illite_img:longname = "Illite refractive index, imag part" ;
		idx_rfr_illite_img:C_format = "%.3g" ;

	float idx_rfr_illite_rl_ee(bnd) ;
		idx_rfr_illite_rl_ee:units = "" ;
		idx_rfr_illite_rl_ee:longname = "Illite refractive index estimated error, real part" ;
		idx_rfr_illite_rl_ee:C_format = "%.4g" ;

	float idx_rfr_illite_img_ee(bnd) ;
		idx_rfr_illite_img_ee:units = "" ;
		idx_rfr_illite_img_ee:longname = "Illite refractive index estimated error, imag part" ;
		idx_rfr_illite_img_ee:C_format = "%.3g" ;

	float idx_rfr_illite_nr(bnd) ;
		idx_rfr_illite_nr:units = "" ;
		idx_rfr_illite_nr:longname = "Illite measured normal reflectance" ;
		idx_rfr_illite_nr:C_format = "%.3g" ;

data:

 bnd_wvn = 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 
    67, 68, 69, 70, 71, 72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 
    85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 
    102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 
    116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 
    130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 
    144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 
    158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 
    172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 
    186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 
    200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 
    214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 
    228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 
    242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 
    256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 
    270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 
    284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 
    298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 
    312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 
    326, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 
    340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 
    354, 355, 356, 357, 358, 359, 360, 361, 362, 363, 364, 365, 366, 367, 
    368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 
    382, 383, 384, 385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395, 
    396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406, 407, 408, 409, 
    410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 
    424, 425, 426, 427, 428, 429, 430, 431, 432, 433, 434, 435, 436, 437, 
    438, 439, 440, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 
    452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 463, 464, 465, 
    466, 467, 468, 469, 470, 471, 472, 473, 474, 475, 476, 477, 478, 479, 
    480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 
    494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 
    508, 509, 510, 511, 512, 513, 514, 515, 516, 517, 518, 519, 520, 521, 
    522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 532, 533, 534, 535, 
    536, 537, 538, 539, 540, 541, 542, 543, 544, 545, 546, 547, 548, 549, 
    550, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563, 
    564, 565, 566, 567, 568, 569, 570, 571, 572, 573, 574, 575, 576, 577, 
    578, 579, 580, 581, 582, 583, 584, 585, 586, 587, 588, 589, 590, 591, 
    592, 593, 594, 595, 596, 597, 598, 599, 600, 601, 602, 603, 604, 605, 
    606, 607, 608, 609, 610, 611, 612, 613, 614, 615, 616, 617, 618, 619, 
    620, 621, 622, 623, 624, 625, 626, 627, 628, 629, 630, 631, 632, 633, 
    634, 635, 636, 637, 638, 639, 640, 641, 642, 643, 644, 645, 646, 647, 
    648, 649, 650, 651, 652, 653, 654, 655, 656, 657, 658, 659, 660, 661, 
    662, 663, 664, 665, 666, 667, 668, 669, 670, 671, 672, 673, 674, 675, 
    676, 677, 678, 679, 680, 681, 682, 683, 684, 685, 686, 687, 688, 689, 
    690, 691, 692, 693, 694, 695, 696, 697, 698, 699, 700, 701, 702, 703, 
    704, 705, 706, 707, 708, 709, 710, 711, 712, 713, 714, 715, 716, 717, 
    718, 719, 720, 721, 722, 723, 724, 725, 726, 727, 728, 729, 730, 731, 
    732, 733, 734, 735, 736, 737, 738, 739, 740, 741, 742, 743, 744, 745, 
    746, 747, 748, 749, 750, 751, 752, 753, 754, 755, 756, 757, 758, 759, 
    760, 761, 762, 763, 764, 765, 766, 767, 768, 769, 770, 771, 772, 773, 
    774, 775, 776, 777, 778, 779, 780, 781, 782, 783, 784, 785, 786, 787, 
    788, 789, 790, 791, 792, 793, 794, 795, 796, 797, 798, 799, 800, 801, 
    802, 803, 804, 805, 806, 807, 808, 809, 810, 811, 812, 813, 814, 815, 
    816, 817, 818, 819, 820, 821, 822, 823, 824, 825, 826, 827, 828, 829, 
    830, 831, 832, 833, 834, 835, 836, 837, 838, 839, 840, 841, 842, 843, 
    844, 845, 846, 847, 848, 849, 850, 851, 852, 853, 854, 855, 856, 857, 
    858, 859, 860, 861, 862, 863, 864, 865, 866, 867, 868, 869, 870, 871, 
    872, 873, 874, 875, 876, 877, 878, 879, 880, 881, 882, 883, 884, 885, 
    886, 887, 888, 889, 890, 891, 892, 893, 894, 895, 896, 897, 898, 899, 
    900, 901, 902, 903, 904, 905, 906, 907, 908, 909, 910, 911, 912, 913, 
    914, 915, 916, 917, 918, 919, 920, 921, 922, 923, 924, 925, 926, 927, 
    928, 929, 930, 931, 932, 933, 934, 935, 936, 937, 938, 939, 940, 941, 
    942, 943, 944, 945, 946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 
    956, 957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 
    970, 971, 972, 973, 974, 975, 976, 977, 978, 979, 980, 981, 982, 983, 
    984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995, 996, 997, 
    998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 
    1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 
    1022, 1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031, 1032, 1033, 
    1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043, 1044, 1045, 
    1046, 1047, 1048, 1049, 1050, 1051, 1052, 1053, 1054, 1055, 1056, 1057, 
    1058, 1059, 1060, 1061, 1062, 1063, 1064, 1065, 1066, 1067, 1068, 1069, 
    1070, 1071, 1072, 1073, 1074, 1075, 1076, 1077, 1078, 1079, 1080, 1081, 
    1082, 1083, 1084, 1085, 1086, 1087, 1088, 1089, 1090, 1091, 1092, 1093, 
    1094, 1095, 1096, 1097, 1098, 1099, 1100, 1101, 1102, 1103, 1104, 1105, 
    1106, 1107, 1108, 1109, 1110, 1111, 1112, 1113, 1114, 1115, 1116, 1117, 
    1118, 1119, 1120, 1121, 1122, 1123, 1124, 1125, 1126, 1127, 1128, 1129, 
    1130, 1131, 1132, 1133, 1134, 1135, 1136, 1137, 1138, 1139, 1140, 1141, 
    1142, 1143, 1144, 1145, 1146, 1147, 1148, 1149, 1150, 1151, 1152, 1153, 
    1154, 1155, 1156, 1157, 1158, 1159, 1160, 1161, 1162, 1163, 1164, 1165, 
    1166, 1167, 1168, 1169, 1170, 1171, 1172, 1173, 1174, 1175, 1176, 1177, 
    1178, 1179, 1180, 1181, 1182, 1183, 1184, 1185, 1186, 1187, 1188, 1189, 
    1190, 1191, 1192, 1193, 1194, 1195, 1196, 1197, 1198, 1199, 1200, 1201, 
    1202, 1203, 1204, 1205, 1206, 1207, 1208, 1209, 1210, 1211, 1212, 1213, 
    1214, 1215, 1216, 1217, 1218, 1219, 1220, 1221, 1222, 1223, 1224, 1225, 
    1226, 1227, 1228, 1229, 1230, 1231, 1232, 1233, 1234, 1235, 1236, 1237, 
    1238, 1239, 1240, 1241, 1242, 1243, 1244, 1245, 1246, 1247, 1248, 1249, 
    1250, 1251, 1252, 1253, 1254, 1255, 1256, 1257, 1258, 1259, 1260, 1261, 
    1262, 1263, 1264, 1265, 1266, 1267, 1268, 1269, 1270, 1271, 1272, 1273, 
    1274, 1275, 1276, 1277, 1278, 1279, 1280, 1281, 1282, 1283, 1284, 1285, 
    1286, 1287, 1288, 1289, 1290, 1291, 1292, 1293, 1294, 1295, 1296, 1297, 
    1298, 1299, 1300, 1301, 1302, 1303, 1304, 1305, 1306, 1307, 1308, 1309, 
    1310, 1311, 1312, 1313, 1314, 1315, 1316, 1317, 1318, 1319, 1320, 1321, 
    1322, 1323, 1324, 1325, 1326, 1327, 1328, 1329, 1330, 1331, 1332, 1333, 
    1334, 1335, 1336, 1337, 1338, 1339, 1340, 1341, 1342, 1343, 1344, 1345, 
    1346, 1347, 1348, 1349, 1350, 1351, 1352, 1353, 1354, 1355, 1356, 1357, 
    1358, 1359, 1360, 1361, 1362, 1363, 1364, 1365, 1366, 1367, 1368, 1369, 
    1370, 1371, 1372, 1373, 1374, 1375, 1376, 1377, 1378, 1379, 1380, 1381, 
    1382, 1383, 1384, 1385, 1386, 1387, 1388, 1389, 1390, 1391, 1392, 1393, 
    1394, 1395, 1396, 1397, 1398, 1399, 1400, 1401, 1402, 1403, 1404, 1405, 
    1406, 1407, 1408, 1409, 1410, 1411, 1412, 1413, 1414, 1415, 1416, 1417, 
    1418, 1419, 1420, 1421, 1422, 1423, 1424, 1425, 1426, 1427, 1428, 1429, 
    1430, 1431, 1432, 1433, 1434, 1435, 1436, 1437, 1438, 1439, 1440, 1441, 
    1442, 1443, 1444, 1445, 1446, 1447, 1448, 1449, 1450, 1451, 1452, 1453, 
    1454, 1455, 1456, 1457, 1458, 1459, 1460, 1461, 1462, 1463, 1464, 1465, 
    1466, 1467, 1468, 1469, 1470, 1471, 1472, 1473, 1474, 1475, 1476, 1477, 
    1478, 1479, 1480, 1481, 1482, 1483, 1484, 1485, 1486, 1487, 1488, 1489, 
    1490, 1491, 1492, 1493, 1494, 1495, 1496, 1497, 1498, 1499, 1500, 1501, 
    1502, 1503, 1504, 1505, 1506, 1507, 1508, 1509, 1510, 1511, 1512, 1513, 
    1514, 1515, 1516, 1517, 1518, 1519, 1520, 1521, 1522, 1523, 1524, 1525, 
    1526, 1527, 1528, 1529, 1530, 1531, 1532, 1533, 1534, 1535, 1536, 1537, 
    1538, 1539, 1540, 1541, 1542, 1543, 1544, 1545, 1546, 1547, 1548, 1549, 
    1550, 1551, 1552, 1553, 1554, 1555, 1556, 1557, 1558, 1559, 1560, 1561, 
    1562, 1563, 1564, 1565, 1566, 1567, 1568, 1569, 1570, 1571, 1572, 1573, 
    1574, 1575, 1576, 1577, 1578, 1579, 1580, 1581, 1582, 1583, 1584, 1585, 
    1586, 1587, 1588, 1589, 1590, 1591, 1592, 1593, 1594, 1595, 1596, 1597, 
    1598, 1599, 1600, 1601, 1602, 1603, 1604, 1605, 1606, 1607, 1608, 1609, 
    1610, 1611, 1612, 1613, 1614, 1615, 1616, 1617, 1618, 1619, 1620, 1621, 
    1622, 1623, 1624, 1625, 1626, 1627, 1628, 1629, 1630, 1631, 1632, 1633, 
    1634, 1635, 1636, 1637, 1638, 1639, 1640, 1641, 1642, 1643, 1644, 1645, 
    1646, 1647, 1648, 1649, 1650, 1651, 1652, 1653, 1654, 1655, 1656, 1657, 
    1658, 1659, 1660, 1661, 1662, 1663, 1664, 1665, 1666, 1667, 1668, 1669, 
    1670, 1671, 1672, 1673, 1674, 1675, 1676, 1677, 1678, 1679, 1680, 1681, 
    1682, 1683, 1684, 1685, 1686, 1687, 1688, 1689, 1690, 1691, 1692, 1693, 
    1694, 1695, 1696, 1697, 1698, 1699, 1700, 1701, 1702, 1703, 1704, 1705, 
    1706, 1707, 1708, 1709, 1710, 1711, 1712, 1713, 1714, 1715, 1716, 1717, 
    1718, 1719, 1720, 1721, 1722, 1723, 1724, 1725, 1726, 1727, 1728, 1729, 
    1730, 1731, 1732, 1733, 1734, 1735, 1736, 1737, 1738, 1739, 1740, 1741, 
    1742, 1743, 1744, 1745, 1746, 1747, 1748, 1749, 1750, 1751, 1752, 1753, 
    1754, 1755, 1756, 1757, 1758, 1759, 1760, 1761, 1762, 1763, 1764, 1765, 
    1766, 1767, 1768, 1769, 1770, 1771, 1772, 1773, 1774, 1775, 1776, 1777, 
    1778, 1779, 1780, 1781, 1782, 1783, 1784, 1785, 1786, 1787, 1788, 1789, 
    1790, 1791, 1792, 1793, 1794, 1795, 1796, 1797, 1798, 1799, 1800, 1801, 
    1802, 1803, 1804, 1805, 1806, 1807, 1808, 1809, 1810, 1811, 1812, 1813, 
    1814, 1815, 1816, 1817, 1818, 1819, 1820, 1821, 1822, 1823, 1824, 1825, 
    1826, 1827, 1828, 1829, 1830, 1831, 1832, 1833, 1834, 1835, 1836, 1837, 
    1838, 1839, 1840, 1841, 1842, 1843, 1844, 1845, 1846, 1847, 1848, 1849, 
    1850, 1851, 1852, 1853, 1854, 1855, 1856, 1857, 1858, 1859, 1860, 1861, 
    1862, 1863, 1864, 1865, 1866, 1867, 1868, 1869, 1870, 1871, 1872, 1873, 
    1874, 1875, 1876, 1877, 1878, 1879, 1880, 1881, 1882, 1883, 1884, 1885, 
    1886, 1887, 1888, 1889, 1890, 1891, 1892, 1893, 1894, 1895, 1896, 1897, 
    1898, 1899, 1900, 1901, 1902, 1903, 1904, 1905, 1906, 1907, 1908, 1909, 
    1910, 1911, 1912, 1913, 1914, 1915, 1916, 1917, 1918, 1919, 1920, 1921, 
    1922, 1923, 1924, 1925, 1926, 1927, 1928, 1929, 1930, 1931, 1932, 1933, 
    1934, 1935, 1936, 1937, 1938, 1939, 1940, 1941, 1942, 1943, 1944, 1945, 
    1946, 1947, 1948, 1949, 1950, 1951, 1952, 1953, 1954, 1955, 1956, 1957, 
    1958, 1959, 1960, 1961, 1962, 1963, 1964, 1965, 1966, 1967, 1968, 1969, 
    1970, 1971, 1972, 1973, 1974, 1975, 1976, 1977, 1978, 1979, 1980, 1981, 
    1982, 1983, 1984, 1985, 1986, 1987, 1988, 1989, 1990, 1991, 1992, 1993, 
    1994, 1995, 1996, 1997, 1998, 1999, 2000, 2001, 2002, 2003, 2004, 2005, 
    2006, 2007, 2008, 2009, 2010, 2011, 2012, 2013, 2014, 2015, 2016, 2017, 
    2018, 2019, 2020, 2021, 2022, 2023, 2024, 2025, 2026, 2027, 2028, 2029, 
    2030, 2031, 2032, 2033, 2034, 2035, 2036, 2037, 2038, 2039, 2040, 2041, 
    2042, 2043, 2044, 2045, 2046, 2047, 2048, 2049, 2050, 2051, 2052, 2053, 
    2054, 2055, 2056, 2057, 2058, 2059, 2060, 2061, 2062, 2063, 2064, 2065, 
    2066, 2067, 2068, 2069, 2070, 2071, 2072, 2073, 2074, 2075, 2076, 2077, 
    2078, 2079, 2080, 2081, 2082, 2083, 2084, 2085, 2086, 2087, 2088, 2089, 
    2090, 2091, 2092, 2093, 2094, 2095, 2096, 2097, 2098, 2099, 2100, 2101, 
    2102, 2103, 2104, 2105, 2106, 2107, 2108, 2109, 2110, 2111, 2112, 2113, 
    2114, 2115, 2116, 2117, 2118, 2119, 2120, 2121, 2122, 2123, 2124, 2125, 
    2126, 2127, 2128, 2129, 2130, 2131, 2132, 2133, 2134, 2135, 2136, 2137, 
    2138, 2139, 2140, 2141, 2142, 2143, 2144, 2145, 2146, 2147, 2148, 2149, 
    2150, 2151, 2152, 2153, 2154, 2155, 2156, 2157, 2158, 2159, 2160, 2161, 
    2162, 2163, 2164, 2165, 2166, 2167, 2168, 2169, 2170, 2171, 2172, 2173, 
    2174, 2175, 2176, 2177, 2178, 2179, 2180, 2181, 2182, 2183, 2184, 2185, 
    2186, 2187, 2188, 2189, 2190, 2191, 2192, 2193, 2194, 2195, 2196, 2197, 
    2198, 2199, 2200, 2201, 2202, 2203, 2204, 2205, 2206, 2207, 2208, 2209, 
    2210, 2211, 2212, 2213, 2214, 2215, 2216, 2217, 2218, 2219, 2220, 2221, 
    2222, 2223, 2224, 2225, 2226, 2227, 2228, 2229, 2230, 2231, 2232, 2233, 
    2234, 2235, 2236, 2237, 2238, 2239, 2240, 2241, 2242, 2243, 2244, 2245, 
    2246, 2247, 2248, 2249, 2250, 2251, 2252, 2253, 2254, 2255, 2256, 2257, 
    2258, 2259, 2260, 2261, 2262, 2263, 2264, 2265, 2266, 2267, 2268, 2269, 
    2270, 2271, 2272, 2273, 2274, 2275, 2276, 2277, 2278, 2279, 2280, 2281, 
    2282, 2283, 2284, 2285, 2286, 2287, 2288, 2289, 2290, 2291, 2292, 2293, 
    2294, 2295, 2296, 2297, 2298, 2299, 2300, 2301, 2302, 2303, 2304, 2305, 
    2306, 2307, 2308, 2309, 2310, 2311, 2312, 2313, 2314, 2315, 2316, 2317, 
    2318, 2319, 2320, 2321, 2322, 2323, 2324, 2325, 2326, 2327, 2328, 2329, 
    2330, 2331, 2332, 2333, 2334, 2335, 2336, 2337, 2338, 2339, 2340, 2341, 
    2342, 2343, 2344, 2345, 2346, 2347, 2348, 2349, 2350, 2351, 2352, 2353, 
    2354, 2355, 2356, 2357, 2358, 2359, 2360, 2361, 2362, 2363, 2364, 2365, 
    2366, 2367, 2368, 2369, 2370, 2371, 2372, 2373, 2374, 2375, 2376, 2377, 
    2378, 2379, 2380, 2381, 2382, 2383, 2384, 2385, 2386, 2387, 2388, 2389, 
    2390, 2391, 2392, 2393, 2394, 2395, 2396, 2397, 2398, 2399, 2400, 2401, 
    2402, 2403, 2404, 2405, 2406, 2407, 2408, 2409, 2410, 2411, 2412, 2413, 
    2414, 2415, 2416, 2417, 2418, 2419, 2420, 2421, 2422, 2423, 2424, 2425, 
    2426, 2427, 2428, 2429, 2430, 2431, 2432, 2433, 2434, 2435, 2436, 2437, 
    2438, 2439, 2440, 2441, 2442, 2443, 2444, 2445, 2446, 2447, 2448, 2449, 
    2450, 2451, 2452, 2453, 2454, 2455, 2456, 2457, 2458, 2459, 2460, 2461, 
    2462, 2463, 2464, 2465, 2466, 2467, 2468, 2469, 2470, 2471, 2472, 2473, 
    2474, 2475, 2476, 2477, 2478, 2479, 2480, 2481, 2482, 2483, 2484, 2485, 
    2486, 2487, 2488, 2489, 2490, 2491, 2492, 2493, 2494, 2495, 2496, 2497, 
    2498, 2499, 2500, 2501, 2502, 2503, 2504, 2505, 2506, 2507, 2508, 2509, 
    2510, 2511, 2512, 2513, 2514, 2515, 2516, 2517, 2518, 2519, 2520, 2521, 
    2522, 2523, 2524, 2525, 2526, 2527, 2528, 2529, 2530, 2531, 2532, 2533, 
    2534, 2535, 2536, 2537, 2538, 2539, 2540, 2541, 2542, 2543, 2544, 2545, 
    2546, 2547, 2548, 2549, 2550, 2551, 2552, 2553, 2554, 2555, 2556, 2557, 
    2558, 2559, 2560, 2561, 2562, 2563, 2564, 2565, 2566, 2567, 2568, 2569, 
    2570, 2571, 2572, 2573, 2574, 2575, 2576, 2577, 2578, 2579, 2580, 2581, 
    2582, 2583, 2584, 2585, 2586, 2587, 2588, 2589, 2590, 2591, 2592, 2593, 
    2594, 2595, 2596, 2597, 2598, 2599, 2600, 2601, 2602, 2603, 2604, 2605, 
    2606, 2607, 2608, 2609, 2610, 2611, 2612, 2613, 2614, 2615, 2616, 2617, 
    2618, 2619, 2620, 2621, 2622, 2623, 2624, 2625, 2626, 2627, 2628, 2629, 
    2630, 2631, 2632, 2633, 2634, 2635, 2636, 2637, 2638, 2639, 2640, 2641, 
    2642, 2643, 2644, 2645, 2646, 2647, 2648, 2649, 2650, 2651, 2652, 2653, 
    2654, 2655, 2656, 2657, 2658, 2659, 2660, 2661, 2662, 2663, 2664, 2665, 
    2666, 2667, 2668, 2669, 2670, 2671, 2672, 2673, 2674, 2675, 2676, 2677, 
    2678, 2679, 2680, 2681, 2682, 2683, 2684, 2685, 2686, 2687, 2688, 2689, 
    2690, 2691, 2692, 2693, 2694, 2695, 2696, 2697, 2698, 2699, 2700, 2701, 
    2702, 2703, 2704, 2705, 2706, 2707, 2708, 2709, 2710, 2711, 2712, 2713, 
    2714, 2715, 2716, 2717, 2718, 2719, 2720, 2721, 2722, 2723, 2724, 2725, 
    2726, 2727, 2728, 2729, 2730, 2731, 2732, 2733, 2734, 2735, 2736, 2737, 
    2738, 2739, 2740, 2741, 2742, 2743, 2744, 2745, 2746, 2747, 2748, 2749, 
    2750, 2751, 2752, 2753, 2754, 2755, 2756, 2757, 2758, 2759, 2760, 2761, 
    2762, 2763, 2764, 2765, 2766, 2767, 2768, 2769, 2770, 2771, 2772, 2773, 
    2774, 2775, 2776, 2777, 2778, 2779, 2780, 2781, 2782, 2783, 2784, 2785, 
    2786, 2787, 2788, 2789, 2790, 2791, 2792, 2793, 2794, 2795, 2796, 2797, 
    2798, 2799, 2800, 2801, 2802, 2803, 2804, 2805, 2806, 2807, 2808, 2809, 
    2810, 2811, 2812, 2813, 2814, 2815, 2816, 2817, 2818, 2819, 2820, 2821, 
    2822, 2823, 2824, 2825, 2826, 2827, 2828, 2829, 2830, 2831, 2832, 2833, 
    2834, 2835, 2836, 2837, 2838, 2839, 2840, 2841, 2842, 2843, 2844, 2845, 
    2846, 2847, 2848, 2849, 2850, 2851, 2852, 2853, 2854, 2855, 2856, 2857, 
    2858, 2859, 2860, 2861, 2862, 2863, 2864, 2865, 2866, 2867, 2868, 2869, 
    2870, 2871, 2872, 2873, 2874, 2875, 2876, 2877, 2878, 2879, 2880, 2881, 
    2882, 2883, 2884, 2885, 2886, 2887, 2888, 2889, 2890, 2891, 2892, 2893, 
    2894, 2895, 2896, 2897, 2898, 2899, 2900, 2901, 2902, 2903, 2904, 2905, 
    2906, 2907, 2908, 2909, 2910, 2911, 2912, 2913, 2914, 2915, 2916, 2917, 
    2918, 2919, 2920, 2921, 2922, 2923, 2924, 2925, 2926, 2927, 2928, 2929, 
    2930, 2931, 2932, 2933, 2934, 2935, 2936, 2937, 2938, 2939, 2940, 2941, 
    2942, 2943, 2944, 2945, 2946, 2947, 2948, 2949, 2950, 2951, 2952, 2953, 
    2954, 2955, 2956, 2957, 2958, 2959, 2960, 2961, 2962, 2963, 2964, 2965, 
    2966, 2967, 2968, 2969, 2970, 2971, 2972, 2973, 2974, 2975, 2976, 2977, 
    2978, 2979, 2980, 2981, 2982, 2983, 2984, 2985, 2986, 2987, 2988, 2989, 
    2990, 2991, 2992, 2993, 2994, 2995, 2996, 2997, 2998, 2999, 3000, 3001, 
    3002, 3003, 3004, 3005, 3006, 3007, 3008, 3009, 3010, 3011, 3012, 3013, 
    3014, 3015, 3016, 3017, 3018, 3019, 3020, 3021, 3022, 3023, 3024, 3025, 
    3026, 3027, 3028, 3029, 3030, 3031, 3032, 3033, 3034, 3035, 3036, 3037, 
    3038, 3039, 3040, 3041, 3042, 3043, 3044, 3045, 3046, 3047, 3048, 3049, 
    3050, 3051, 3052, 3053, 3054, 3055, 3056, 3057, 3058, 3059, 3060, 3061, 
    3062, 3063, 3064, 3065, 3066, 3067, 3068, 3069, 3070, 3071, 3072, 3073, 
    3074, 3075, 3076, 3077, 3078, 3079, 3080, 3081, 3082, 3083, 3084, 3085, 
    3086, 3087, 3088, 3089, 3090, 3091, 3092, 3093, 3094, 3095, 3096, 3097, 
    3098, 3099, 3100, 3101, 3102, 3103, 3104, 3105, 3106, 3107, 3108, 3109, 
    3110, 3111, 3112, 3113, 3114, 3115, 3116, 3117, 3118, 3119, 3120, 3121, 
    3122, 3123, 3124, 3125, 3126, 3127, 3128, 3129, 3130, 3131, 3132, 3133, 
    3134, 3135, 3136, 3137, 3138, 3139, 3140, 3141, 3142, 3143, 3144, 3145, 
    3146, 3147, 3148, 3149, 3150, 3151, 3152, 3153, 3154, 3155, 3156, 3157, 
    3158, 3159, 3160, 3161, 3162, 3163, 3164, 3165, 3166, 3167, 3168, 3169, 
    3170, 3171, 3172, 3173, 3174, 3175, 3176, 3177, 3178, 3179, 3180, 3181, 
    3182, 3183, 3184, 3185, 3186, 3187, 3188, 3189, 3190, 3191, 3192, 3193, 
    3194, 3195, 3196, 3197, 3198, 3199, 3200, 3201, 3202, 3203, 3204, 3205, 
    3206, 3207, 3208, 3209, 3210, 3211, 3212, 3213, 3214, 3215, 3216, 3217, 
    3218, 3219, 3220, 3221, 3222, 3223, 3224, 3225, 3226, 3227, 3228, 3229, 
    3230, 3231, 3232, 3233, 3234, 3235, 3236, 3237, 3238, 3239, 3240, 3241, 
    3242, 3243, 3244, 3245, 3246, 3247, 3248, 3249, 3250, 3251, 3252, 3253, 
    3254, 3255, 3256, 3257, 3258, 3259, 3260, 3261, 3262, 3263, 3264, 3265, 
    3266, 3267, 3268, 3269, 3270, 3271, 3272, 3273, 3274, 3275, 3276, 3277, 
    3278, 3279, 3280, 3281, 3282, 3283, 3284, 3285, 3286, 3287, 3288, 3289, 
    3290, 3291, 3292, 3293, 3294, 3295, 3296, 3297, 3298, 3299, 3300, 3301, 
    3302, 3303, 3304, 3305, 3306, 3307, 3308, 3309, 3310, 3311, 3312, 3313, 
    3314, 3315, 3316, 3317, 3318, 3319, 3320, 3321, 3322, 3323, 3324, 3325, 
    3326, 3327, 3328, 3329, 3330, 3331, 3332, 3333, 3334, 3335, 3336, 3337, 
    3338, 3339, 3340, 3341, 3342, 3343, 3344, 3345, 3346, 3347, 3348, 3349, 
    3350, 3351, 3352, 3353, 3354, 3355, 3356, 3357, 3358, 3359, 3360, 3361, 
    3362, 3363, 3364, 3365, 3366, 3367, 3368, 3369, 3370, 3371, 3372, 3373, 
    3374, 3375, 3376, 3377, 3378, 3379, 3380, 3381, 3382, 3383, 3384, 3385, 
    3386, 3387, 3388, 3389, 3390, 3391, 3392, 3393, 3394, 3395, 3396, 3397, 
    3398, 3399, 3400, 3401, 3402, 3403, 3404, 3405, 3406, 3407, 3408, 3409, 
    3410, 3411, 3412, 3413, 3414, 3415, 3416, 3417, 3418, 3419, 3420, 3421, 
    3422, 3423, 3424, 3425, 3426, 3427, 3428, 3429, 3430, 3431, 3432, 3433, 
    3434, 3435, 3436, 3437, 3438, 3439, 3440, 3441, 3442, 3443, 3444, 3445, 
    3446, 3447, 3448, 3449, 3450, 3451, 3452, 3453, 3454, 3455, 3456, 3457, 
    3458, 3459, 3460, 3461, 3462, 3463, 3464, 3465, 3466, 3467, 3468, 3469, 
    3470, 3471, 3472, 3473, 3474, 3475, 3476, 3477, 3478, 3479, 3480, 3481, 
    3482, 3483, 3484, 3485, 3486, 3487, 3488, 3489, 3490, 3491, 3492, 3493, 
    3494, 3495, 3496, 3497, 3498, 3499, 3500, 3501, 3502, 3503, 3504, 3505, 
    3506, 3507, 3508, 3509, 3510, 3511, 3512, 3513, 3514, 3515, 3516, 3517, 
    3518, 3519, 3520, 3521, 3522, 3523, 3524, 3525, 3526, 3527, 3528, 3529, 
    3530, 3531, 3532, 3533, 3534, 3535, 3536, 3537, 3538, 3539, 3540, 3541, 
    3542, 3543, 3544, 3545, 3546, 3547, 3548, 3549, 3550, 3551, 3552, 3553, 
    3554, 3555, 3556, 3557, 3558, 3559, 3560, 3561, 3562, 3563, 3564, 3565, 
    3566, 3567, 3568, 3569, 3570, 3571, 3572, 3573, 3574, 3575, 3576, 3577, 
    3578, 3579, 3580, 3581, 3582, 3583, 3584, 3585, 3586, 3587, 3588, 3589, 
    3590, 3591, 3592, 3593, 3594, 3595, 3596, 3597, 3598, 3599, 3600, 3601, 
    3602, 3603, 3604, 3605, 3606, 3607, 3608, 3609, 3610, 3611, 3612, 3613, 
    3614, 3615, 3616, 3617, 3618, 3619, 3620, 3621, 3622, 3623, 3624, 3625, 
    3626, 3627, 3628, 3629, 3630, 3631, 3632, 3633, 3634, 3635, 3636, 3637, 
    3638, 3639, 3640, 3641, 3642, 3643, 3644, 3645, 3646, 3647, 3648, 3649, 
    3650, 3651, 3652, 3653, 3654, 3655, 3656, 3657, 3658, 3659, 3660, 3661, 
    3662, 3663, 3664, 3665, 3666, 3667, 3668, 3669, 3670, 3671, 3672, 3673, 
    3674, 3675, 3676, 3677, 3678, 3679, 3680, 3681, 3682, 3683, 3684, 3685, 
    3686, 3687, 3688, 3689, 3690, 3691, 3692, 3693, 3694, 3695, 3696, 3697, 
    3698, 3699, 3700, 3701, 3702, 3703, 3704, 3705, 3706, 3707, 3708, 3709, 
    3710, 3711, 3712, 3713, 3714, 3715, 3716, 3717, 3718, 3719, 3720, 3721, 
    3722, 3723, 3724, 3725, 3726, 3727, 3728, 3729, 3730, 3731, 3732, 3733, 
    3734, 3735, 3736, 3737, 3738, 3739, 3740, 3741, 3742, 3743, 3744, 3745, 
    3746, 3747, 3748, 3749, 3750, 3751, 3752, 3753, 3754, 3755, 3756, 3757, 
    3758, 3759, 3760, 3761, 3762, 3763, 3764, 3765, 3766, 3767, 3768, 3769, 
    3770, 3771, 3772, 3773, 3774, 3775, 3776, 3777, 3778, 3779, 3780, 3781, 
    3782, 3783, 3784, 3785, 3786, 3787, 3788, 3789, 3790, 3791, 3792, 3793, 
    3794, 3795, 3796, 3797, 3798, 3799, 3800, 3801, 3802, 3803, 3804, 3805, 
    3806, 3807, 3808, 3809, 3810, 3811, 3812, 3813, 3814, 3815, 3816, 3817, 
    3818, 3819, 3820, 3821, 3822, 3823, 3824, 3825, 3826, 3827, 3828, 3829, 
    3830, 3831, 3832, 3833, 3834, 3835, 3836, 3837, 3838, 3839, 3840, 3841, 
    3842, 3843, 3844, 3845, 3846, 3847, 3848, 3849, 3850, 3851, 3852, 3853, 
    3854, 3855, 3856, 3857, 3858, 3859, 3860, 3861, 3862, 3863, 3864, 3865, 
    3866, 3867, 3868, 3869, 3870, 3871, 3872, 3873, 3874, 3875, 3876, 3877, 
    3878, 3879, 3880, 3881, 3882, 3883, 3884, 3885, 3886, 3887, 3888, 3889, 
    3890, 3891, 3892, 3893, 3894, 3895, 3896, 3897, 3898, 3899, 3900, 3901, 
    3902, 3903, 3904, 3905, 3906, 3907, 3908, 3909, 3910, 3911, 3912, 3913, 
    3914, 3915, 3916, 3917, 3918, 3919, 3920, 3921, 3922, 3923, 3924, 3925, 
    3926, 3927, 3928, 3929, 3930, 3931, 3932, 3933, 3934, 3935, 3936, 3937, 
    3938, 3939, 3940, 3941, 3942, 3943, 3944, 3945, 3946, 3947, 3948, 3949, 
    3950, 3951, 3952, 3953, 3954, 3955, 3956, 3957, 3958, 3959, 3960, 3961, 
    3962, 3963, 3964, 3965, 3966, 3967, 3968, 3969, 3970, 3971, 3972, 3973, 
    3974, 3975, 3976, 3977, 3978, 3979, 3980, 3981, 3982, 3983, 3984, 3985, 
    3986, 3987, 3988, 3989, 3990, 3991, 3992, 3993, 3994, 3995, 3996, 3997, 
    3998, 3999, 4000 ;

 bnd = 200, 196.08, 192.31, 188.68, 185.19, 181.82, 178.57, 175.44, 
    172.41, 169.49, 166.67, 163.93, 161.29, 158.73, 156.25, 153.85, 151.52, 
    149.25, 147.06, 144.93, 142.86, 140.85, 138.89, 136.99, 135.14, 133.33, 
    131.58, 129.87, 128.21, 126.58, 125, 123.46, 121.95, 120.48, 119.05, 
    117.65, 116.28, 114.94, 113.64, 112.36, 111.11, 109.89, 108.7, 107.53, 
    106.38, 105.26, 104.17, 103.09, 102.04, 101.01, 100, 99.01, 98.039, 
    97.087, 96.154, 95.238, 94.34, 93.458, 92.593, 91.743, 90.909, 90.09, 
    89.286, 88.496, 87.719, 86.956, 86.207, 85.47, 84.746, 84.034, 83.333, 
    82.645, 81.967, 81.301, 80.645, 80, 79.365, 78.74, 78.125, 77.519, 
    76.923, 76.336, 75.758, 75.188, 74.627, 74.074, 73.529, 72.993, 72.464, 
    71.942, 71.429, 70.922, 70.423, 69.93, 69.444, 68.965, 68.493, 68.027, 
    67.568, 67.114, 66.667, 66.225, 65.789, 65.359, 64.935, 64.516, 64.103, 
    63.694, 63.291, 62.893, 62.5, 62.112, 61.728, 61.35, 60.976, 60.606, 
    60.241, 59.88, 59.524, 59.172, 58.824, 58.479, 58.139, 57.804, 57.471, 
    57.143, 56.818, 56.497, 56.18, 55.866, 55.556, 55.249, 54.945, 54.645, 
    54.348, 54.054, 53.763, 53.476, 53.192, 52.91, 52.632, 52.356, 52.083, 
    51.813, 51.546, 51.282, 51.02, 50.761, 50.505, 50.251, 50, 49.751, 
    49.505, 49.261, 49.02, 48.78, 48.544, 48.309, 48.077, 47.847, 47.619, 
    47.393, 47.17, 46.948, 46.729, 46.512, 46.296, 46.083, 45.872, 45.662, 
    45.454, 45.249, 45.045, 44.843, 44.643, 44.444, 44.248, 44.053, 43.86, 
    43.668, 43.478, 43.29, 43.103, 42.918, 42.735, 42.553, 42.373, 42.194, 
    42.017, 41.841, 41.667, 41.494, 41.322, 41.152, 40.984, 40.816, 40.65, 
    40.486, 40.323, 40.161, 40, 39.841, 39.682, 39.526, 39.37, 39.216, 
    39.062, 38.91, 38.76, 38.61, 38.461, 38.314, 38.168, 38.023, 37.879, 
    37.736, 37.594, 37.453, 37.313, 37.175, 37.037, 36.9, 36.765, 36.63, 
    36.496, 36.364, 36.232, 36.101, 35.971, 35.842, 35.714, 35.587, 35.461, 
    35.336, 35.211, 35.088, 34.965, 34.843, 34.722, 34.602, 34.483, 34.364, 
    34.247, 34.13, 34.014, 33.898, 33.784, 33.67, 33.557, 33.445, 33.333, 
    33.223, 33.113, 33.003, 32.895, 32.787, 32.68, 32.573, 32.467, 32.362, 
    32.258, 32.154, 32.051, 31.949, 31.847, 31.746, 31.646, 31.546, 31.447, 
    31.348, 31.25, 31.153, 31.056, 30.96, 30.864, 30.769, 30.675, 30.581, 
    30.488, 30.395, 30.303, 30.212, 30.121, 30.03, 29.94, 29.851, 29.762, 
    29.674, 29.586, 29.499, 29.412, 29.326, 29.24, 29.154, 29.07, 28.986, 
    28.902, 28.818, 28.736, 28.653, 28.571, 28.49, 28.409, 28.329, 28.249, 
    28.169, 28.09, 28.011, 27.933, 27.855, 27.778, 27.701, 27.624, 27.548, 
    27.472, 27.397, 27.322, 27.248, 27.174, 27.1, 27.027, 26.954, 26.882, 
    26.81, 26.738, 26.667, 26.596, 26.525, 26.455, 26.385, 26.316, 26.247, 
    26.178, 26.11, 26.042, 25.974, 25.907, 25.84, 25.773, 25.707, 25.641, 
    25.575, 25.51, 25.445, 25.381, 25.316, 25.253, 25.189, 25.126, 25.063, 
    25, 24.938, 24.876, 24.814, 24.753, 24.691, 24.631, 24.57, 24.51, 24.45, 
    24.39, 24.331, 24.272, 24.213, 24.155, 24.096, 24.038, 23.981, 23.923, 
    23.866, 23.809, 23.753, 23.697, 23.641, 23.585, 23.529, 23.474, 23.419, 
    23.365, 23.31, 23.256, 23.202, 23.148, 23.095, 23.042, 22.989, 22.936, 
    22.883, 22.831, 22.779, 22.727, 22.676, 22.624, 22.573, 22.522, 22.472, 
    22.421, 22.371, 22.321, 22.272, 22.222, 22.173, 22.124, 22.075, 22.026, 
    21.978, 21.93, 21.882, 21.834, 21.787, 21.739, 21.692, 21.645, 21.598, 
    21.552, 21.505, 21.459, 21.413, 21.368, 21.322, 21.277, 21.231, 21.186, 
    21.142, 21.097, 21.053, 21.008, 20.964, 20.92, 20.877, 20.833, 20.79, 
    20.747, 20.704, 20.661, 20.619, 20.576, 20.534, 20.492, 20.45, 20.408, 
    20.367, 20.325, 20.284, 20.243, 20.202, 20.161, 20.121, 20.08, 20.04, 20, 
    19.96, 19.92, 19.881, 19.841, 19.802, 19.763, 19.724, 19.685, 19.646, 
    19.608, 19.569, 19.531, 19.493, 19.455, 19.417, 19.38, 19.342, 19.305, 
    19.268, 19.231, 19.194, 19.157, 19.121, 19.084, 19.048, 19.011, 18.975, 
    18.939, 18.904, 18.868, 18.832, 18.797, 18.762, 18.727, 18.692, 18.657, 
    18.622, 18.587, 18.553, 18.518, 18.484, 18.45, 18.416, 18.382, 18.349, 
    18.315, 18.281, 18.248, 18.215, 18.182, 18.149, 18.116, 18.083, 18.051, 
    18.018, 17.986, 17.953, 17.921, 17.889, 17.857, 17.825, 17.794, 17.762, 
    17.73, 17.699, 17.668, 17.637, 17.606, 17.575, 17.544, 17.513, 17.483, 
    17.452, 17.422, 17.391, 17.361, 17.331, 17.301, 17.271, 17.241, 17.212, 
    17.182, 17.153, 17.123, 17.094, 17.065, 17.036, 17.007, 16.978, 16.949, 
    16.92, 16.892, 16.863, 16.835, 16.807, 16.778, 16.75, 16.722, 16.694, 
    16.667, 16.639, 16.611, 16.584, 16.556, 16.529, 16.502, 16.475, 16.447, 
    16.42, 16.393, 16.367, 16.34, 16.313, 16.287, 16.26, 16.234, 16.208, 
    16.181, 16.155, 16.129, 16.103, 16.077, 16.051, 16.026, 16, 15.974, 
    15.949, 15.924, 15.898, 15.873, 15.848, 15.823, 15.798, 15.773, 15.748, 
    15.723, 15.699, 15.674, 15.649, 15.625, 15.601, 15.576, 15.552, 15.528, 
    15.504, 15.48, 15.456, 15.432, 15.408, 15.385, 15.361, 15.337, 15.314, 
    15.29, 15.267, 15.244, 15.221, 15.198, 15.175, 15.151, 15.129, 15.106, 
    15.083, 15.06, 15.038, 15.015, 14.993, 14.97, 14.948, 14.925, 14.903, 
    14.881, 14.859, 14.837, 14.815, 14.793, 14.771, 14.749, 14.727, 14.706, 
    14.684, 14.663, 14.641, 14.62, 14.599, 14.577, 14.556, 14.535, 14.514, 
    14.493, 14.472, 14.451, 14.43, 14.409, 14.389, 14.368, 14.347, 14.327, 
    14.306, 14.286, 14.265, 14.245, 14.225, 14.205, 14.184, 14.164, 14.144, 
    14.124, 14.104, 14.085, 14.065, 14.045, 14.025, 14.006, 13.986, 13.967, 
    13.947, 13.928, 13.908, 13.889, 13.87, 13.85, 13.831, 13.812, 13.793, 
    13.774, 13.755, 13.736, 13.717, 13.699, 13.68, 13.661, 13.643, 13.624, 
    13.605, 13.587, 13.568, 13.55, 13.532, 13.514, 13.495, 13.477, 13.459, 
    13.441, 13.423, 13.405, 13.387, 13.369, 13.351, 13.333, 13.316, 13.298, 
    13.28, 13.263, 13.245, 13.227, 13.21, 13.193, 13.175, 13.158, 13.141, 
    13.123, 13.106, 13.089, 13.072, 13.055, 13.038, 13.021, 13.004, 12.987, 
    12.97, 12.953, 12.937, 12.92, 12.903, 12.887, 12.87, 12.854, 12.837, 
    12.821, 12.804, 12.788, 12.771, 12.755, 12.739, 12.723, 12.707, 12.69, 
    12.674, 12.658, 12.642, 12.626, 12.61, 12.594, 12.579, 12.563, 12.547, 
    12.531, 12.516, 12.5, 12.484, 12.469, 12.453, 12.438, 12.422, 12.407, 
    12.392, 12.376, 12.361, 12.346, 12.33, 12.315, 12.3, 12.285, 12.27, 
    12.255, 12.24, 12.225, 12.21, 12.195, 12.18, 12.165, 12.151, 12.136, 
    12.121, 12.106, 12.092, 12.077, 12.063, 12.048, 12.034, 12.019, 12.005, 
    11.99, 11.976, 11.962, 11.947, 11.933, 11.919, 11.905, 11.891, 11.877, 
    11.862, 11.848, 11.834, 11.82, 11.806, 11.792, 11.779, 11.765, 11.751, 
    11.737, 11.723, 11.71, 11.696, 11.682, 11.669, 11.655, 11.641, 11.628, 
    11.614, 11.601, 11.587, 11.574, 11.561, 11.547, 11.534, 11.521, 11.507, 
    11.494, 11.481, 11.468, 11.455, 11.442, 11.429, 11.415, 11.403, 11.389, 
    11.377, 11.364, 11.351, 11.338, 11.325, 11.312, 11.299, 11.287, 11.274, 
    11.261, 11.249, 11.236, 11.223, 11.211, 11.198, 11.186, 11.173, 11.161, 
    11.148, 11.136, 11.123, 11.111, 11.099, 11.087, 11.074, 11.062, 11.05, 
    11.038, 11.025, 11.013, 11.001, 10.989, 10.977, 10.965, 10.953, 10.941, 
    10.929, 10.917, 10.905, 10.893, 10.881, 10.87, 10.858, 10.846, 10.834, 
    10.823, 10.811, 10.799, 10.788, 10.776, 10.764, 10.753, 10.741, 10.73, 
    10.718, 10.707, 10.695, 10.684, 10.672, 10.661, 10.65, 10.638, 10.627, 
    10.616, 10.604, 10.593, 10.582, 10.571, 10.56, 10.549, 10.537, 10.526, 
    10.515, 10.504, 10.493, 10.482, 10.471, 10.46, 10.449, 10.438, 10.427, 
    10.417, 10.406, 10.395, 10.384, 10.373, 10.363, 10.352, 10.341, 10.331, 
    10.32, 10.309, 10.299, 10.288, 10.278, 10.267, 10.256, 10.246, 10.235, 
    10.225, 10.215, 10.204, 10.194, 10.183, 10.173, 10.163, 10.152, 10.142, 
    10.132, 10.122, 10.111, 10.101, 10.091, 10.081, 10.071, 10.06, 10.05, 
    10.04, 10.03, 10.02, 10.01, 10, 9.99, 9.98, 9.9701, 9.9602, 9.9502, 
    9.9404, 9.9305, 9.9206, 9.9108, 9.901, 9.8912, 9.8814, 9.8717, 9.8619, 
    9.8522, 9.8425, 9.8328, 9.8232, 9.8135, 9.8039, 9.7943, 9.7847, 9.7752, 
    9.7656, 9.7561, 9.7466, 9.7371, 9.7276, 9.7182, 9.7087, 9.6993, 9.6899, 
    9.6805, 9.6712, 9.6618, 9.6525, 9.6432, 9.6339, 9.6246, 9.6154, 9.6061, 
    9.5969, 9.5877, 9.5785, 9.5694, 9.5602, 9.5511, 9.542, 9.5329, 9.5238, 
    9.5147, 9.5057, 9.4967, 9.4877, 9.4787, 9.4697, 9.4607, 9.4518, 9.4429, 
    9.434, 9.4251, 9.4162, 9.4073, 9.3985, 9.3897, 9.3809, 9.3721, 9.3633, 
    9.3545, 9.3458, 9.3371, 9.3284, 9.3197, 9.311, 9.3023, 9.2937, 9.2851, 
    9.2764, 9.2678, 9.2593, 9.2507, 9.2421, 9.2336, 9.2251, 9.2166, 9.2081, 
    9.1996, 9.1912, 9.1827, 9.1743, 9.1659, 9.1575, 9.1491, 9.1408, 9.1324, 
    9.1241, 9.1158, 9.1075, 9.0992, 9.0909, 9.0827, 9.0744, 9.0662, 9.058, 
    9.0498, 9.0416, 9.0334, 9.0253, 9.0171, 9.009, 9.0009, 8.9928, 8.9847, 
    8.9767, 8.9686, 8.9606, 8.9526, 8.9445, 8.9366, 8.9286, 8.9206, 8.9127, 
    8.9047, 8.8968, 8.8889, 8.881, 8.8731, 8.8652, 8.8574, 8.8496, 8.8417, 
    8.8339, 8.8261, 8.8183, 8.8106, 8.8028, 8.7951, 8.7873, 8.7796, 8.7719, 
    8.7642, 8.7566, 8.7489, 8.7413, 8.7336, 8.726, 8.7184, 8.7108, 8.7032, 
    8.6957, 8.6881, 8.6806, 8.673, 8.6655, 8.658, 8.6505, 8.643, 8.6356, 
    8.6281, 8.6207, 8.6133, 8.6059, 8.5985, 8.5911, 8.5837, 8.5763, 8.569, 
    8.5616, 8.5543, 8.547, 8.5397, 8.5324, 8.5251, 8.5179, 8.5106, 8.5034, 
    8.4962, 8.489, 8.4818, 8.4746, 8.4674, 8.4602, 8.4531, 8.4459, 8.4388, 
    8.4317, 8.4246, 8.4175, 8.4104, 8.4034, 8.3963, 8.3893, 8.3822, 8.3752, 
    8.3682, 8.3612, 8.3542, 8.3472, 8.3403, 8.3333, 8.3264, 8.3195, 8.3126, 
    8.3056, 8.2988, 8.2919, 8.285, 8.2781, 8.2713, 8.2645, 8.2576, 8.2508, 
    8.244, 8.2372, 8.2305, 8.2237, 8.2169, 8.2102, 8.2034, 8.1967, 8.19, 
    8.1833, 8.1766, 8.1699, 8.1633, 8.1566, 8.15, 8.1433, 8.1367, 8.1301, 
    8.1235, 8.1169, 8.1103, 8.1037, 8.0972, 8.0906, 8.0841, 8.0775, 8.071, 
    8.0645, 8.058, 8.0515, 8.0451, 8.0386, 8.0321, 8.0257, 8.0192, 8.0128, 
    8.0064, 8, 7.9936, 7.9872, 7.9808, 7.9745, 7.9681, 7.9618, 7.9554, 
    7.9491, 7.9428, 7.9365, 7.9302, 7.9239, 7.9177, 7.9114, 7.9051, 7.8989, 
    7.8927, 7.8864, 7.8802, 7.874, 7.8678, 7.8616, 7.8555, 7.8493, 7.8431, 
    7.837, 7.8309, 7.8247, 7.8186, 7.8125, 7.8064, 7.8003, 7.7942, 7.7882, 
    7.7821, 7.776, 7.77, 7.764, 7.758, 7.7519, 7.7459, 7.7399, 7.734, 7.728, 
    7.722, 7.716, 7.7101, 7.7042, 7.6982, 7.6923, 7.6864, 7.6805, 7.6746, 
    7.6687, 7.6628, 7.657, 7.6511, 7.6453, 7.6394, 7.6336, 7.6278, 7.622, 
    7.6161, 7.6104, 7.6046, 7.5988, 7.593, 7.5873, 7.5815, 7.5758, 7.57, 
    7.5643, 7.5586, 7.5529, 7.5472, 7.5415, 7.5358, 7.5301, 7.5245, 7.5188, 
    7.5131, 7.5075, 7.5019, 7.4963, 7.4906, 7.485, 7.4794, 7.4738, 7.4683, 
    7.4627, 7.4571, 7.4516, 7.446, 7.4405, 7.4349, 7.4294, 7.4239, 7.4184, 
    7.4129, 7.4074, 7.4019, 7.3964, 7.391, 7.3855, 7.3801, 7.3746, 7.3692, 
    7.3638, 7.3584, 7.3529, 7.3475, 7.3421, 7.3368, 7.3314, 7.326, 7.3206, 
    7.3153, 7.3099, 7.3046, 7.2993, 7.2939, 7.2886, 7.2833, 7.278, 7.2727, 
    7.2674, 7.2622, 7.2569, 7.2516, 7.2464, 7.2411, 7.2359, 7.2307, 7.2254, 
    7.2202, 7.215, 7.2098, 7.2046, 7.1994, 7.1942, 7.1891, 7.1839, 7.1788, 
    7.1736, 7.1685, 7.1633, 7.1582, 7.1531, 7.148, 7.1429, 7.1378, 7.1327, 
    7.1276, 7.1225, 7.1174, 7.1124, 7.1073, 7.1023, 7.0972, 7.0922, 7.0872, 
    7.0822, 7.0771, 7.0721, 7.0671, 7.0621, 7.0572, 7.0522, 7.0472, 7.0423, 
    7.0373, 7.0323, 7.0274, 7.0225, 7.0175, 7.0126, 7.0077, 7.0028, 6.9979, 
    6.993, 6.9881, 6.9832, 6.9784, 6.9735, 6.9686, 6.9638, 6.9589, 6.9541, 
    6.9493, 6.9444, 6.9396, 6.9348, 6.93, 6.9252, 6.9204, 6.9156, 6.9109, 
    6.9061, 6.9013, 6.8966, 6.8918, 6.8871, 6.8823, 6.8776, 6.8729, 6.8681, 
    6.8634, 6.8587, 6.854, 6.8493, 6.8446, 6.8399, 6.8353, 6.8306, 6.8259, 
    6.8213, 6.8166, 6.812, 6.8074, 6.8027, 6.7981, 6.7935, 6.7889, 6.7843, 
    6.7797, 6.7751, 6.7705, 6.7659, 6.7613, 6.7568, 6.7522, 6.7476, 6.7431, 
    6.7385, 6.734, 6.7295, 6.7249, 6.7204, 6.7159, 6.7114, 6.7069, 6.7024, 
    6.6979, 6.6934, 6.689, 6.6845, 6.68, 6.6756, 6.6711, 6.6667, 6.6622, 
    6.6578, 6.6534, 6.6489, 6.6445, 6.6401, 6.6357, 6.6313, 6.6269, 6.6225, 
    6.6181, 6.6138, 6.6094, 6.605, 6.6007, 6.5963, 6.592, 6.5876, 6.5833, 
    6.5789, 6.5746, 6.5703, 6.566, 6.5617, 6.5574, 6.5531, 6.5488, 6.5445, 
    6.5402, 6.5359, 6.5317, 6.5274, 6.5232, 6.5189, 6.5147, 6.5104, 6.5062, 
    6.502, 6.4977, 6.4935, 6.4893, 6.4851, 6.4809, 6.4767, 6.4725, 6.4683, 
    6.4641, 6.4599, 6.4558, 6.4516, 6.4475, 6.4433, 6.4392, 6.435, 6.4309, 
    6.4267, 6.4226, 6.4185, 6.4144, 6.4103, 6.4061, 6.402, 6.398, 6.3939, 
    6.3898, 6.3857, 6.3816, 6.3776, 6.3735, 6.3694, 6.3654, 6.3613, 6.3573, 
    6.3532, 6.3492, 6.3452, 6.3412, 6.3371, 6.3331, 6.3291, 6.3251, 6.3211, 
    6.3171, 6.3131, 6.3091, 6.3052, 6.3012, 6.2972, 6.2933, 6.2893, 6.2854, 
    6.2814, 6.2775, 6.2735, 6.2696, 6.2657, 6.2617, 6.2578, 6.2539, 6.25, 
    6.2461, 6.2422, 6.2383, 6.2344, 6.2305, 6.2267, 6.2228, 6.2189, 6.215, 
    6.2112, 6.2073, 6.2035, 6.1996, 6.1958, 6.192, 6.1881, 6.1843, 6.1805, 
    6.1767, 6.1728, 6.169, 6.1652, 6.1614, 6.1576, 6.1538, 6.1501, 6.1463, 
    6.1425, 6.1387, 6.135, 6.1312, 6.1275, 6.1237, 6.12, 6.1162, 6.1125, 
    6.1087, 6.105, 6.1013, 6.0976, 6.0938, 6.0901, 6.0864, 6.0827, 6.079, 
    6.0753, 6.0716, 6.068, 6.0643, 6.0606, 6.0569, 6.0533, 6.0496, 6.0459, 
    6.0423, 6.0386, 6.035, 6.0314, 6.0277, 6.0241, 6.0205, 6.0168, 6.0132, 
    6.0096, 6.006, 6.0024, 5.9988, 5.9952, 5.9916, 5.988, 5.9844, 5.9809, 
    5.9773, 5.9737, 5.9701, 5.9666, 5.963, 5.9595, 5.9559, 5.9524, 5.9488, 
    5.9453, 5.9418, 5.9382, 5.9347, 5.9312, 5.9277, 5.9242, 5.9207, 5.9172, 
    5.9137, 5.9102, 5.9067, 5.9032, 5.8997, 5.8962, 5.8928, 5.8893, 5.8858, 
    5.8824, 5.8789, 5.8754, 5.872, 5.8685, 5.8651, 5.8617, 5.8582, 5.8548, 
    5.8514, 5.848, 5.8445, 5.8411, 5.8377, 5.8343, 5.8309, 5.8275, 5.8241, 
    5.8207, 5.8173, 5.814, 5.8106, 5.8072, 5.8038, 5.8005, 5.7971, 5.7937, 
    5.7904, 5.787, 5.7837, 5.7803, 5.777, 5.7737, 5.7703, 5.767, 5.7637, 
    5.7604, 5.7571, 5.7537, 5.7504, 5.7471, 5.7438, 5.7405, 5.7372, 5.7339, 
    5.7307, 5.7274, 5.7241, 5.7208, 5.7176, 5.7143, 5.711, 5.7078, 5.7045, 
    5.7013, 5.698, 5.6948, 5.6915, 5.6883, 5.685, 5.6818, 5.6786, 5.6754, 
    5.6721, 5.6689, 5.6657, 5.6625, 5.6593, 5.6561, 5.6529, 5.6497, 5.6465, 
    5.6433, 5.6402, 5.637, 5.6338, 5.6306, 5.6275, 5.6243, 5.6211, 5.618, 
    5.6148, 5.6117, 5.6085, 5.6054, 5.6022, 5.5991, 5.596, 5.5928, 5.5897, 
    5.5866, 5.5835, 5.5804, 5.5772, 5.5741, 5.571, 5.5679, 5.5648, 5.5617, 
    5.5586, 5.5556, 5.5525, 5.5494, 5.5463, 5.5432, 5.5402, 5.5371, 5.534, 
    5.531, 5.5279, 5.5249, 5.5218, 5.5188, 5.5157, 5.5127, 5.5096, 5.5066, 
    5.5036, 5.5006, 5.4975, 5.4945, 5.4915, 5.4885, 5.4855, 5.4825, 5.4795, 
    5.4765, 5.4735, 5.4705, 5.4675, 5.4645, 5.4615, 5.4585, 5.4555, 5.4526, 
    5.4496, 5.4466, 5.4437, 5.4407, 5.4377, 5.4348, 5.4318, 5.4289, 5.4259, 
    5.423, 5.4201, 5.4171, 5.4142, 5.4113, 5.4083, 5.4054, 5.4025, 5.3996, 
    5.3967, 5.3937, 5.3908, 5.3879, 5.385, 5.3821, 5.3792, 5.3763, 5.3735, 
    5.3706, 5.3677, 5.3648, 5.3619, 5.3591, 5.3562, 5.3533, 5.3505, 5.3476, 
    5.3447, 5.3419, 5.339, 5.3362, 5.3333, 5.3305, 5.3277, 5.3248, 5.322, 
    5.3191, 5.3163, 5.3135, 5.3107, 5.3079, 5.305, 5.3022, 5.2994, 5.2966, 
    5.2938, 5.291, 5.2882, 5.2854, 5.2826, 5.2798, 5.277, 5.2743, 5.2715, 
    5.2687, 5.2659, 5.2632, 5.2604, 5.2576, 5.2549, 5.2521, 5.2493, 5.2466, 
    5.2438, 5.2411, 5.2383, 5.2356, 5.2329, 5.2301, 5.2274, 5.2247, 5.2219, 
    5.2192, 5.2165, 5.2138, 5.211, 5.2083, 5.2056, 5.2029, 5.2002, 5.1975, 
    5.1948, 5.1921, 5.1894, 5.1867, 5.184, 5.1813, 5.1787, 5.176, 5.1733, 
    5.1706, 5.168, 5.1653, 5.1626, 5.16, 5.1573, 5.1546, 5.152, 5.1493, 
    5.1467, 5.144, 5.1414, 5.1387, 5.1361, 5.1335, 5.1308, 5.1282, 5.1256, 
    5.123, 5.1203, 5.1177, 5.1151, 5.1125, 5.1099, 5.1073, 5.1046, 5.102, 
    5.0994, 5.0968, 5.0942, 5.0916, 5.0891, 5.0865, 5.0839, 5.0813, 5.0787, 
    5.0761, 5.0736, 5.071, 5.0684, 5.0659, 5.0633, 5.0607, 5.0582, 5.0556, 
    5.0531, 5.0505, 5.048, 5.0454, 5.0429, 5.0403, 5.0378, 5.0352, 5.0327, 
    5.0302, 5.0277, 5.0251, 5.0226, 5.0201, 5.0176, 5.015, 5.0125, 5.01, 
    5.0075, 5.005, 5.0025, 5, 4.9975, 4.995, 4.9925, 4.99, 4.9875, 4.985, 
    4.9826, 4.9801, 4.9776, 4.9751, 4.9727, 4.9702, 4.9677, 4.9652, 4.9628, 
    4.9603, 4.9579, 4.9554, 4.9529, 4.9505, 4.948, 4.9456, 4.9432, 4.9407, 
    4.9383, 4.9358, 4.9334, 4.931, 4.9285, 4.9261, 4.9237, 4.9213, 4.9188, 
    4.9164, 4.914, 4.9116, 4.9092, 4.9068, 4.9044, 4.902, 4.8996, 4.8972, 
    4.8948, 4.8924, 4.89, 4.8876, 4.8852, 4.8828, 4.8804, 4.878, 4.8757, 
    4.8733, 4.8709, 4.8685, 4.8662, 4.8638, 4.8614, 4.8591, 4.8567, 4.8544, 
    4.852, 4.8497, 4.8473, 4.845, 4.8426, 4.8403, 4.8379, 4.8356, 4.8333, 
    4.8309, 4.8286, 4.8263, 4.8239, 4.8216, 4.8193, 4.817, 4.8146, 4.8123, 
    4.81, 4.8077, 4.8054, 4.8031, 4.8008, 4.7985, 4.7962, 4.7939, 4.7916, 
    4.7893, 4.787, 4.7847, 4.7824, 4.7801, 4.7778, 4.7755, 4.7733, 4.771, 
    4.7687, 4.7664, 4.7642, 4.7619, 4.7596, 4.7574, 4.7551, 4.7529, 4.7506, 
    4.7483, 4.7461, 4.7438, 4.7416, 4.7393, 4.7371, 4.7348, 4.7326, 4.7304, 
    4.7281, 4.7259, 4.7237, 4.7214, 4.7192, 4.717, 4.7148, 4.7125, 4.7103, 
    4.7081, 4.7059, 4.7037, 4.7015, 4.6992, 4.697, 4.6948, 4.6926, 4.6904, 
    4.6882, 4.686, 4.6838, 4.6816, 4.6795, 4.6773, 4.6751, 4.6729, 4.6707, 
    4.6685, 4.6664, 4.6642, 4.662, 4.6598, 4.6577, 4.6555, 4.6533, 4.6512, 
    4.649, 4.6468, 4.6447, 4.6425, 4.6404, 4.6382, 4.6361, 4.6339, 4.6318, 
    4.6296, 4.6275, 4.6253, 4.6232, 4.6211, 4.6189, 4.6168, 4.6147, 4.6125, 
    4.6104, 4.6083, 4.6062, 4.6041, 4.6019, 4.5998, 4.5977, 4.5956, 4.5935, 
    4.5914, 4.5893, 4.5872, 4.5851, 4.583, 4.5809, 4.5788, 4.5767, 4.5746, 
    4.5725, 4.5704, 4.5683, 4.5662, 4.5641, 4.562, 4.56, 4.5579, 4.5558, 
    4.5537, 4.5517, 4.5496, 4.5475, 4.5455, 4.5434, 4.5413, 4.5393, 4.5372, 
    4.5351, 4.5331, 4.531, 4.529, 4.5269, 4.5249, 4.5228, 4.5208, 4.5188, 
    4.5167, 4.5147, 4.5126, 4.5106, 4.5086, 4.5065, 4.5045, 4.5025, 4.5005, 
    4.4984, 4.4964, 4.4944, 4.4924, 4.4903, 4.4883, 4.4863, 4.4843, 4.4823, 
    4.4803, 4.4783, 4.4763, 4.4743, 4.4723, 4.4703, 4.4683, 4.4663, 4.4643, 
    4.4623, 4.4603, 4.4583, 4.4563, 4.4543, 4.4524, 4.4504, 4.4484, 4.4464, 
    4.4444, 4.4425, 4.4405, 4.4385, 4.4366, 4.4346, 4.4326, 4.4307, 4.4287, 
    4.4267, 4.4248, 4.4228, 4.4209, 4.4189, 4.417, 4.415, 4.4131, 4.4111, 
    4.4092, 4.4072, 4.4053, 4.4033, 4.4014, 4.3995, 4.3975, 4.3956, 4.3937, 
    4.3917, 4.3898, 4.3879, 4.386, 4.384, 4.3821, 4.3802, 4.3783, 4.3764, 
    4.3745, 4.3725, 4.3706, 4.3687, 4.3668, 4.3649, 4.363, 4.3611, 4.3592, 
    4.3573, 4.3554, 4.3535, 4.3516, 4.3497, 4.3478, 4.3459, 4.344, 4.3422, 
    4.3403, 4.3384, 4.3365, 4.3346, 4.3328, 4.3309, 4.329, 4.3271, 4.3253, 
    4.3234, 4.3215, 4.3197, 4.3178, 4.3159, 4.3141, 4.3122, 4.3103, 4.3085, 
    4.3066, 4.3048, 4.3029, 4.3011, 4.2992, 4.2974, 4.2955, 4.2937, 4.2918, 
    4.29, 4.2882, 4.2863, 4.2845, 4.2827, 4.2808, 4.279, 4.2772, 4.2753, 
    4.2735, 4.2717, 4.2699, 4.268, 4.2662, 4.2644, 4.2626, 4.2608, 4.2589, 
    4.2571, 4.2553, 4.2535, 4.2517, 4.2499, 4.2481, 4.2463, 4.2445, 4.2427, 
    4.2409, 4.2391, 4.2373, 4.2355, 4.2337, 4.2319, 4.2301, 4.2283, 4.2265, 
    4.2248, 4.223, 4.2212, 4.2194, 4.2176, 4.2159, 4.2141, 4.2123, 4.2105, 
    4.2088, 4.207, 4.2052, 4.2034, 4.2017, 4.1999, 4.1982, 4.1964, 4.1946, 
    4.1929, 4.1911, 4.1894, 4.1876, 4.1859, 4.1841, 4.1824, 4.1806, 4.1789, 
    4.1771, 4.1754, 4.1736, 4.1719, 4.1701, 4.1684, 4.1667, 4.1649, 4.1632, 
    4.1615, 4.1597, 4.158, 4.1563, 4.1545, 4.1528, 4.1511, 4.1494, 4.1477, 
    4.1459, 4.1442, 4.1425, 4.1408, 4.1391, 4.1374, 4.1356, 4.1339, 4.1322, 
    4.1305, 4.1288, 4.1271, 4.1254, 4.1237, 4.122, 4.1203, 4.1186, 4.1169, 
    4.1152, 4.1135, 4.1118, 4.1102, 4.1085, 4.1068, 4.1051, 4.1034, 4.1017, 
    4.1, 4.0984, 4.0967, 4.095, 4.0933, 4.0917, 4.09, 4.0883, 4.0866, 4.085, 
    4.0833, 4.0816, 4.08, 4.0783, 4.0766, 4.075, 4.0733, 4.0717, 4.07, 
    4.0683, 4.0667, 4.065, 4.0634, 4.0617, 4.0601, 4.0584, 4.0568, 4.0552, 
    4.0535, 4.0519, 4.0502, 4.0486, 4.0469, 4.0453, 4.0437, 4.042, 4.0404, 
    4.0388, 4.0371, 4.0355, 4.0339, 4.0323, 4.0306, 4.029, 4.0274, 4.0258, 
    4.0241, 4.0225, 4.0209, 4.0193, 4.0177, 4.0161, 4.0145, 4.0128, 4.0112, 
    4.0096, 4.008, 4.0064, 4.0048, 4.0032, 4.0016, 4, 3.9984, 3.9968, 3.9952, 
    3.9936, 3.992, 3.9904, 3.9888, 3.9872, 3.9857, 3.9841, 3.9825, 3.9809, 
    3.9793, 3.9777, 3.9761, 3.9746, 3.973, 3.9714, 3.9698, 3.9683, 3.9667, 
    3.9651, 3.9635, 3.962, 3.9604, 3.9588, 3.9573, 3.9557, 3.9541, 3.9526, 
    3.951, 3.9494, 3.9479, 3.9463, 3.9448, 3.9432, 3.9417, 3.9401, 3.9386, 
    3.937, 3.9355, 3.9339, 3.9324, 3.9308, 3.9293, 3.9277, 3.9262, 3.9246, 
    3.9231, 3.9216, 3.92, 3.9185, 3.917, 3.9154, 3.9139, 3.9124, 3.9108, 
    3.9093, 3.9078, 3.9063, 3.9047, 3.9032, 3.9017, 3.9002, 3.8986, 3.8971, 
    3.8956, 3.8941, 3.8926, 3.8911, 3.8895, 3.888, 3.8865, 3.885, 3.8835, 
    3.882, 3.8805, 3.879, 3.8775, 3.876, 3.8745, 3.873, 3.8715, 3.87, 3.8685, 
    3.867, 3.8655, 3.864, 3.8625, 3.861, 3.8595, 3.858, 3.8565, 3.8551, 
    3.8536, 3.8521, 3.8506, 3.8491, 3.8476, 3.8462, 3.8447, 3.8432, 3.8417, 
    3.8402, 3.8388, 3.8373, 3.8358, 3.8344, 3.8329, 3.8314, 3.83, 3.8285, 
    3.827, 3.8256, 3.8241, 3.8226, 3.8212, 3.8197, 3.8183, 3.8168, 3.8153, 
    3.8139, 3.8124, 3.811, 3.8095, 3.8081, 3.8066, 3.8052, 3.8037, 3.8023, 
    3.8008, 3.7994, 3.7979, 3.7965, 3.7951, 3.7936, 3.7922, 3.7908, 3.7893, 
    3.7879, 3.7864, 3.785, 3.7836, 3.7821, 3.7807, 3.7793, 3.7779, 3.7764, 
    3.775, 3.7736, 3.7722, 3.7707, 3.7693, 3.7679, 3.7665, 3.7651, 3.7636, 
    3.7622, 3.7608, 3.7594, 3.758, 3.7566, 3.7552, 3.7538, 3.7523, 3.7509, 
    3.7495, 3.7481, 3.7467, 3.7453, 3.7439, 3.7425, 3.7411, 3.7397, 3.7383, 
    3.7369, 3.7355, 3.7341, 3.7327, 3.7313, 3.73, 3.7286, 3.7272, 3.7258, 
    3.7244, 3.723, 3.7216, 3.7202, 3.7189, 3.7175, 3.7161, 3.7147, 3.7133, 
    3.712, 3.7106, 3.7092, 3.7078, 3.7064, 3.7051, 3.7037, 3.7023, 3.701, 
    3.6996, 3.6982, 3.6969, 3.6955, 3.6941, 3.6928, 3.6914, 3.69, 3.6887, 
    3.6873, 3.686, 3.6846, 3.6832, 3.6819, 3.6805, 3.6792, 3.6778, 3.6765, 
    3.6751, 3.6738, 3.6724, 3.6711, 3.6697, 3.6684, 3.667, 3.6657, 3.6643, 
    3.663, 3.6617, 3.6603, 3.659, 3.6576, 3.6563, 3.655, 3.6536, 3.6523, 
    3.651, 3.6496, 3.6483, 3.647, 3.6456, 3.6443, 3.643, 3.6417, 3.6403, 
    3.639, 3.6377, 3.6364, 3.635, 3.6337, 3.6324, 3.6311, 3.6298, 3.6284, 
    3.6271, 3.6258, 3.6245, 3.6232, 3.6219, 3.6206, 3.6193, 3.6179, 3.6166, 
    3.6153, 3.614, 3.6127, 3.6114, 3.6101, 3.6088, 3.6075, 3.6062, 3.6049, 
    3.6036, 3.6023, 3.601, 3.5997, 3.5984, 3.5971, 3.5958, 3.5945, 3.5932, 
    3.592, 3.5907, 3.5894, 3.5881, 3.5868, 3.5855, 3.5842, 3.5829, 3.5817, 
    3.5804, 3.5791, 3.5778, 3.5765, 3.5753, 3.574, 3.5727, 3.5714, 3.5702, 
    3.5689, 3.5676, 3.5663, 3.5651, 3.5638, 3.5625, 3.5613, 3.56, 3.5587, 
    3.5575, 3.5562, 3.5549, 3.5537, 3.5524, 3.5511, 3.5499, 3.5486, 3.5474, 
    3.5461, 3.5448, 3.5436, 3.5423, 3.5411, 3.5398, 3.5386, 3.5373, 3.5361, 
    3.5348, 3.5336, 3.5323, 3.5311, 3.5298, 3.5286, 3.5273, 3.5261, 3.5249, 
    3.5236, 3.5224, 3.5211, 3.5199, 3.5186, 3.5174, 3.5162, 3.5149, 3.5137, 
    3.5125, 3.5112, 3.51, 3.5088, 3.5075, 3.5063, 3.5051, 3.5039, 3.5026, 
    3.5014, 3.5002, 3.499, 3.4977, 3.4965, 3.4953, 3.4941, 3.4928, 3.4916, 
    3.4904, 3.4892, 3.488, 3.4868, 3.4855, 3.4843, 3.4831, 3.4819, 3.4807, 
    3.4795, 3.4783, 3.4771, 3.4758, 3.4746, 3.4734, 3.4722, 3.471, 3.4698, 
    3.4686, 3.4674, 3.4662, 3.465, 3.4638, 3.4626, 3.4614, 3.4602, 3.459, 
    3.4578, 3.4566, 3.4554, 3.4542, 3.453, 3.4518, 3.4507, 3.4495, 3.4483, 
    3.4471, 3.4459, 3.4447, 3.4435, 3.4423, 3.4412, 3.44, 3.4388, 3.4376, 
    3.4364, 3.4352, 3.4341, 3.4329, 3.4317, 3.4305, 3.4294, 3.4282, 3.427, 
    3.4258, 3.4247, 3.4235, 3.4223, 3.4211, 3.42, 3.4188, 3.4176, 3.4165, 
    3.4153, 3.4141, 3.413, 3.4118, 3.4106, 3.4095, 3.4083, 3.4072, 3.406, 
    3.4048, 3.4037, 3.4025, 3.4014, 3.4002, 3.399, 3.3979, 3.3967, 3.3956, 
    3.3944, 3.3933, 3.3921, 3.391, 3.3898, 3.3887, 3.3875, 3.3864, 3.3852, 
    3.3841, 3.3829, 3.3818, 3.3807, 3.3795, 3.3784, 3.3772, 3.3761, 3.375, 
    3.3738, 3.3727, 3.3715, 3.3704, 3.3693, 3.3681, 3.367, 3.3659, 3.3647, 
    3.3636, 3.3625, 3.3613, 3.3602, 3.3591, 3.358, 3.3568, 3.3557, 3.3546, 
    3.3535, 3.3523, 3.3512, 3.3501, 3.349, 3.3478, 3.3467, 3.3456, 3.3445, 
    3.3434, 3.3422, 3.3411, 3.34, 3.3389, 3.3378, 3.3367, 3.3356, 3.3344, 
    3.3333, 3.3322, 3.3311, 3.33, 3.3289, 3.3278, 3.3267, 3.3256, 3.3245, 
    3.3234, 3.3223, 3.3212, 3.3201, 3.319, 3.3179, 3.3167, 3.3156, 3.3146, 
    3.3135, 3.3124, 3.3113, 3.3102, 3.3091, 3.308, 3.3069, 3.3058, 3.3047, 
    3.3036, 3.3025, 3.3014, 3.3003, 3.2992, 3.2982, 3.2971, 3.296, 3.2949, 
    3.2938, 3.2927, 3.2916, 3.2906, 3.2895, 3.2884, 3.2873, 3.2862, 3.2852, 
    3.2841, 3.283, 3.2819, 3.2808, 3.2798, 3.2787, 3.2776, 3.2765, 3.2755, 
    3.2744, 3.2733, 3.2723, 3.2712, 3.2701, 3.269, 3.268, 3.2669, 3.2658, 
    3.2648, 3.2637, 3.2626, 3.2616, 3.2605, 3.2595, 3.2584, 3.2573, 3.2563, 
    3.2552, 3.2541, 3.2531, 3.252, 3.251, 3.2499, 3.2489, 3.2478, 3.2468, 
    3.2457, 3.2446, 3.2436, 3.2425, 3.2415, 3.2404, 3.2394, 3.2383, 3.2373, 
    3.2362, 3.2352, 3.2342, 3.2331, 3.2321, 3.231, 3.23, 3.2289, 3.2279, 
    3.2268, 3.2258, 3.2248, 3.2237, 3.2227, 3.2216, 3.2206, 3.2196, 3.2185, 
    3.2175, 3.2165, 3.2154, 3.2144, 3.2134, 3.2123, 3.2113, 3.2103, 3.2092, 
    3.2082, 3.2072, 3.2062, 3.2051, 3.2041, 3.2031, 3.202, 3.201, 3.2, 3.199, 
    3.198, 3.1969, 3.1959, 3.1949, 3.1939, 3.1928, 3.1918, 3.1908, 3.1898, 
    3.1888, 3.1878, 3.1867, 3.1857, 3.1847, 3.1837, 3.1827, 3.1817, 3.1807, 
    3.1797, 3.1786, 3.1776, 3.1766, 3.1756, 3.1746, 3.1736, 3.1726, 3.1716, 
    3.1706, 3.1696, 3.1686, 3.1676, 3.1666, 3.1656, 3.1646, 3.1636, 3.1626, 
    3.1616, 3.1606, 3.1596, 3.1586, 3.1576, 3.1566, 3.1556, 3.1546, 3.1536, 
    3.1526, 3.1516, 3.1506, 3.1496, 3.1486, 3.1476, 3.1466, 3.1456, 3.1447, 
    3.1437, 3.1427, 3.1417, 3.1407, 3.1397, 3.1387, 3.1377, 3.1368, 3.1358, 
    3.1348, 3.1338, 3.1328, 3.1319, 3.1309, 3.1299, 3.1289, 3.1279, 3.127, 
    3.126, 3.125, 3.124, 3.123, 3.1221, 3.1211, 3.1201, 3.1192, 3.1182, 
    3.1172, 3.1162, 3.1153, 3.1143, 3.1133, 3.1124, 3.1114, 3.1104, 3.1095, 
    3.1085, 3.1075, 3.1066, 3.1056, 3.1046, 3.1037, 3.1027, 3.1017, 3.1008, 
    3.0998, 3.0989, 3.0979, 3.0969, 3.096, 3.095, 3.0941, 3.0931, 3.0921, 
    3.0912, 3.0902, 3.0893, 3.0883, 3.0874, 3.0864, 3.0855, 3.0845, 3.0836, 
    3.0826, 3.0817, 3.0807, 3.0798, 3.0788, 3.0779, 3.0769, 3.076, 3.075, 
    3.0741, 3.0731, 3.0722, 3.0713, 3.0703, 3.0694, 3.0684, 3.0675, 3.0665, 
    3.0656, 3.0647, 3.0637, 3.0628, 3.0618, 3.0609, 3.06, 3.059, 3.0581, 
    3.0572, 3.0562, 3.0553, 3.0544, 3.0534, 3.0525, 3.0516, 3.0506, 3.0497, 
    3.0488, 3.0479, 3.0469, 3.046, 3.0451, 3.0441, 3.0432, 3.0423, 3.0414, 
    3.0404, 3.0395, 3.0386, 3.0377, 3.0367, 3.0358, 3.0349, 3.034, 3.0331, 
    3.0321, 3.0312, 3.0303, 3.0294, 3.0285, 3.0276, 3.0266, 3.0257, 3.0248, 
    3.0239, 3.023, 3.0221, 3.0211, 3.0202, 3.0193, 3.0184, 3.0175, 3.0166, 
    3.0157, 3.0148, 3.0139, 3.013, 3.012, 3.0111, 3.0102, 3.0093, 3.0084, 
    3.0075, 3.0066, 3.0057, 3.0048, 3.0039, 3.003, 3.0021, 3.0012, 3.0003, 
    2.9994, 2.9985, 2.9976, 2.9967, 2.9958, 2.9949, 2.994, 2.9931, 2.9922, 
    2.9913, 2.9904, 2.9895, 2.9886, 2.9878, 2.9869, 2.986, 2.9851, 2.9842, 
    2.9833, 2.9824, 2.9815, 2.9806, 2.9797, 2.9789, 2.978, 2.9771, 2.9762, 
    2.9753, 2.9744, 2.9735, 2.9727, 2.9718, 2.9709, 2.97, 2.9691, 2.9682, 
    2.9674, 2.9665, 2.9656, 2.9647, 2.9638, 2.963, 2.9621, 2.9612, 2.9603, 
    2.9595, 2.9586, 2.9577, 2.9568, 2.956, 2.9551, 2.9542, 2.9533, 2.9525, 
    2.9516, 2.9507, 2.9499, 2.949, 2.9481, 2.9472, 2.9464, 2.9455, 2.9446, 
    2.9438, 2.9429, 2.942, 2.9412, 2.9403, 2.9394, 2.9386, 2.9377, 2.9369, 
    2.936, 2.9351, 2.9343, 2.9334, 2.9326, 2.9317, 2.9308, 2.93, 2.9291, 
    2.9283, 2.9274, 2.9265, 2.9257, 2.9248, 2.924, 2.9231, 2.9223, 2.9214, 
    2.9206, 2.9197, 2.9189, 2.918, 2.9172, 2.9163, 2.9155, 2.9146, 2.9138, 
    2.9129, 2.9121, 2.9112, 2.9104, 2.9095, 2.9087, 2.9078, 2.907, 2.9061, 
    2.9053, 2.9044, 2.9036, 2.9028, 2.9019, 2.9011, 2.9002, 2.8994, 2.8986, 
    2.8977, 2.8969, 2.896, 2.8952, 2.8944, 2.8935, 2.8927, 2.8918, 2.891, 
    2.8902, 2.8893, 2.8885, 2.8877, 2.8868, 2.886, 2.8852, 2.8843, 2.8835, 
    2.8827, 2.8818, 2.881, 2.8802, 2.8794, 2.8785, 2.8777, 2.8769, 2.876, 
    2.8752, 2.8744, 2.8736, 2.8727, 2.8719, 2.8711, 2.8703, 2.8694, 2.8686, 
    2.8678, 2.867, 2.8662, 2.8653, 2.8645, 2.8637, 2.8629, 2.862, 2.8612, 
    2.8604, 2.8596, 2.8588, 2.858, 2.8571, 2.8563, 2.8555, 2.8547, 2.8539, 
    2.8531, 2.8523, 2.8514, 2.8506, 2.8498, 2.849, 2.8482, 2.8474, 2.8466, 
    2.8458, 2.845, 2.8441, 2.8433, 2.8425, 2.8417, 2.8409, 2.8401, 2.8393, 
    2.8385, 2.8377, 2.8369, 2.8361, 2.8353, 2.8345, 2.8337, 2.8329, 2.8321, 
    2.8313, 2.8305, 2.8297, 2.8289, 2.8281, 2.8273, 2.8265, 2.8257, 2.8249, 
    2.8241, 2.8233, 2.8225, 2.8217, 2.8209, 2.8201, 2.8193, 2.8185, 2.8177, 
    2.8169, 2.8161, 2.8153, 2.8145, 2.8137, 2.8129, 2.8121, 2.8114, 2.8106, 
    2.8098, 2.809, 2.8082, 2.8074, 2.8066, 2.8058, 2.805, 2.8043, 2.8035, 
    2.8027, 2.8019, 2.8011, 2.8003, 2.7996, 2.7988, 2.798, 2.7972, 2.7964, 
    2.7956, 2.7949, 2.7941, 2.7933, 2.7925, 2.7917, 2.791, 2.7902, 2.7894, 
    2.7886, 2.7878, 2.7871, 2.7863, 2.7855, 2.7847, 2.784, 2.7832, 2.7824, 
    2.7816, 2.7809, 2.7801, 2.7793, 2.7785, 2.7778, 2.777, 2.7762, 2.7755, 
    2.7747, 2.7739, 2.7732, 2.7724, 2.7716, 2.7709, 2.7701, 2.7693, 2.7685, 
    2.7678, 2.767, 2.7663, 2.7655, 2.7647, 2.764, 2.7632, 2.7624, 2.7617, 
    2.7609, 2.7601, 2.7594, 2.7586, 2.7579, 2.7571, 2.7563, 2.7556, 2.7548, 
    2.7541, 2.7533, 2.7525, 2.7518, 2.751, 2.7503, 2.7495, 2.7488, 2.748, 
    2.7473, 2.7465, 2.7457, 2.745, 2.7442, 2.7435, 2.7427, 2.742, 2.7412, 
    2.7405, 2.7397, 2.739, 2.7382, 2.7375, 2.7367, 2.736, 2.7352, 2.7345, 
    2.7337, 2.733, 2.7322, 2.7315, 2.7307, 2.73, 2.7293, 2.7285, 2.7278, 
    2.727, 2.7263, 2.7255, 2.7248, 2.7241, 2.7233, 2.7226, 2.7218, 2.7211, 
    2.7203, 2.7196, 2.7189, 2.7181, 2.7174, 2.7167, 2.7159, 2.7152, 2.7144, 
    2.7137, 2.713, 2.7122, 2.7115, 2.7108, 2.71, 2.7093, 2.7086, 2.7078, 
    2.7071, 2.7064, 2.7056, 2.7049, 2.7042, 2.7034, 2.7027, 2.702, 2.7012, 
    2.7005, 2.6998, 2.6991, 2.6983, 2.6976, 2.6969, 2.6961, 2.6954, 2.6947, 
    2.694, 2.6932, 2.6925, 2.6918, 2.6911, 2.6903, 2.6896, 2.6889, 2.6882, 
    2.6874, 2.6867, 2.686, 2.6853, 2.6846, 2.6838, 2.6831, 2.6824, 2.6817, 
    2.681, 2.6802, 2.6795, 2.6788, 2.6781, 2.6774, 2.6767, 2.6759, 2.6752, 
    2.6745, 2.6738, 2.6731, 2.6724, 2.6717, 2.6709, 2.6702, 2.6695, 2.6688, 
    2.6681, 2.6674, 2.6667, 2.666, 2.6652, 2.6645, 2.6638, 2.6631, 2.6624, 
    2.6617, 2.661, 2.6603, 2.6596, 2.6589, 2.6582, 2.6575, 2.6567, 2.656, 
    2.6553, 2.6546, 2.6539, 2.6532, 2.6525, 2.6518, 2.6511, 2.6504, 2.6497, 
    2.649, 2.6483, 2.6476, 2.6469, 2.6462, 2.6455, 2.6448, 2.6441, 2.6434, 
    2.6427, 2.642, 2.6413, 2.6406, 2.6399, 2.6392, 2.6385, 2.6378, 2.6371, 
    2.6364, 2.6357, 2.635, 2.6344, 2.6337, 2.633, 2.6323, 2.6316, 2.6309, 
    2.6302, 2.6295, 2.6288, 2.6281, 2.6274, 2.6267, 2.6261, 2.6254, 2.6247, 
    2.624, 2.6233, 2.6226, 2.6219, 2.6212, 2.6205, 2.6199, 2.6192, 2.6185, 
    2.6178, 2.6171, 2.6164, 2.6157, 2.6151, 2.6144, 2.6137, 2.613, 2.6123, 
    2.6116, 2.611, 2.6103, 2.6096, 2.6089, 2.6082, 2.6076, 2.6069, 2.6062, 
    2.6055, 2.6048, 2.6042, 2.6035, 2.6028, 2.6021, 2.6015, 2.6008, 2.6001, 
    2.5994, 2.5988, 2.5981, 2.5974, 2.5967, 2.5961, 2.5954, 2.5947, 2.594, 
    2.5934, 2.5927, 2.592, 2.5913, 2.5907, 2.59, 2.5893, 2.5887, 2.588, 
    2.5873, 2.5867, 2.586, 2.5853, 2.5846, 2.584, 2.5833, 2.5826, 2.582, 
    2.5813, 2.5806, 2.58, 2.5793, 2.5786, 2.578, 2.5773, 2.5767, 2.576, 
    2.5753, 2.5747, 2.574, 2.5733, 2.5727, 2.572, 2.5714, 2.5707, 2.57, 
    2.5694, 2.5687, 2.5681, 2.5674, 2.5667, 2.5661, 2.5654, 2.5648, 2.5641, 
    2.5634, 2.5628, 2.5621, 2.5615, 2.5608, 2.5602, 2.5595, 2.5589, 2.5582, 
    2.5575, 2.5569, 2.5562, 2.5556, 2.5549, 2.5543, 2.5536, 2.553, 2.5523, 
    2.5517, 2.551, 2.5504, 2.5497, 2.5491, 2.5484, 2.5478, 2.5471, 2.5465, 
    2.5458, 2.5452, 2.5445, 2.5439, 2.5432, 2.5426, 2.5419, 2.5413, 2.5407, 
    2.54, 2.5394, 2.5387, 2.5381, 2.5374, 2.5368, 2.5361, 2.5355, 2.5349, 
    2.5342, 2.5336, 2.5329, 2.5323, 2.5316, 2.531, 2.5304, 2.5297, 2.5291, 
    2.5284, 2.5278, 2.5272, 2.5265, 2.5259, 2.5253, 2.5246, 2.524, 2.5233, 
    2.5227, 2.5221, 2.5214, 2.5208, 2.5202, 2.5195, 2.5189, 2.5183, 2.5176, 
    2.517, 2.5164, 2.5157, 2.5151, 2.5145, 2.5138, 2.5132, 2.5126, 2.5119, 
    2.5113, 2.5107, 2.51, 2.5094, 2.5088, 2.5082, 2.5075, 2.5069, 2.5063, 
    2.5056, 2.505, 2.5044, 2.5038, 2.5031, 2.5025, 2.5019, 2.5013, 2.5006, 2.5 ;

 idx_rfr_illite_rl = 2.188, 2.19, 2.191, 2.194, 2.196, 2.199, 2.202, 2.206, 
    2.21, 2.214, 2.217, 2.221, 2.224, 2.228, 2.233, 2.239, 2.245, 2.252, 
    2.259, 2.267, 2.274, 2.282, 2.289, 2.296, 2.303, 2.312, 2.322, 2.33, 
    2.339, 2.346, 2.352, 2.355, 2.357, 2.356, 2.353, 2.348, 2.343, 2.338, 
    2.331, 2.322, 2.313, 2.303, 2.291, 2.28, 2.268, 2.254, 2.24, 2.227, 
    2.214, 2.201, 2.187, 2.174, 2.159, 2.145, 2.13, 2.114, 2.097, 2.078, 
    2.06, 2.043, 2.028, 2.015, 2.005, 1.999, 1.996, 1.995, 1.996, 1.998, 2, 
    2.001, 2.002, 2.002, 2.003, 2.002, 2.003, 2.003, 2.002, 2.001, 1.999, 
    1.997, 1.993, 1.99, 1.986, 1.982, 1.978, 1.975, 1.973, 1.971, 1.971, 
    1.972, 1.972, 1.974, 1.975, 1.976, 1.978, 1.979, 1.98, 1.982, 1.983, 
    1.985, 1.986, 1.988, 1.99, 1.992, 1.993, 1.994, 1.995, 1.995, 1.995, 
    1.995, 1.995, 1.994, 1.995, 1.996, 1.997, 2, 2.003, 2.006, 2.01, 2.014, 
    2.018, 2.022, 2.025, 2.029, 2.032, 2.034, 2.037, 2.039, 2.04, 2.041, 
    2.041, 2.041, 2.039, 2.037, 2.033, 2.029, 2.024, 2.02, 2.015, 2.012, 
    2.009, 2.006, 2.004, 2.002, 2.001, 2, 1.999, 1.999, 1.999, 1.999, 2.001, 
    2.003, 2.006, 2.009, 2.012, 2.015, 2.019, 2.023, 2.027, 2.031, 2.034, 
    2.036, 2.039, 2.041, 2.042, 2.044, 2.045, 2.047, 2.05, 2.053, 2.057, 
    2.06, 2.063, 2.065, 2.067, 2.07, 2.072, 2.074, 2.077, 2.081, 2.085, 
    2.088, 2.091, 2.094, 2.097, 2.101, 2.104, 2.107, 2.111, 2.115, 2.12, 
    2.124, 2.128, 2.131, 2.134, 2.135, 2.136, 2.136, 2.136, 2.134, 2.132, 
    2.129, 2.126, 2.122, 2.117, 2.112, 2.106, 2.1, 2.093, 2.086, 2.079, 
    2.072, 2.065, 2.057, 2.051, 2.044, 2.039, 2.034, 2.03, 2.028, 2.027, 
    2.026, 2.028, 2.03, 2.032, 2.036, 2.04, 2.044, 2.049, 2.054, 2.058, 
    2.062, 2.066, 2.07, 2.074, 2.078, 2.081, 2.085, 2.088, 2.092, 2.096, 
    2.099, 2.102, 2.106, 2.11, 2.114, 2.118, 2.122, 2.126, 2.13, 2.134, 
    2.138, 2.143, 2.147, 2.15, 2.154, 2.158, 2.161, 2.164, 2.168, 2.171, 
    2.174, 2.177, 2.18, 2.182, 2.185, 2.188, 2.19, 2.192, 2.195, 2.197, 
    2.199, 2.201, 2.204, 2.207, 2.21, 2.213, 2.216, 2.219, 2.223, 2.226, 
    2.23, 2.233, 2.237, 2.242, 2.247, 2.252, 2.257, 2.263, 2.269, 2.274, 
    2.28, 2.284, 2.289, 2.292, 2.295, 2.296, 2.296, 2.296, 2.294, 2.291, 
    2.288, 2.284, 2.28, 2.276, 2.271, 2.267, 2.264, 2.261, 2.258, 2.256, 
    2.254, 2.252, 2.249, 2.245, 2.24, 2.234, 2.227, 2.217, 2.207, 2.196, 
    2.185, 2.174, 2.164, 2.156, 2.15, 2.146, 2.145, 2.147, 2.152, 2.159, 
    2.17, 2.182, 2.197, 2.214, 2.231, 2.248, 2.264, 2.278, 2.29, 2.298, 
    2.302, 2.301, 2.298, 2.291, 2.282, 2.271, 2.262, 2.253, 2.248, 2.245, 
    2.246, 2.252, 2.261, 2.273, 2.289, 2.306, 2.324, 2.342, 2.36, 2.376, 
    2.39, 2.402, 2.411, 2.417, 2.421, 2.423, 2.423, 2.422, 2.418, 2.414, 
    2.408, 2.401, 2.392, 2.383, 2.373, 2.363, 2.352, 2.341, 2.331, 2.322, 
    2.313, 2.306, 2.3, 2.296, 2.294, 2.293, 2.295, 2.298, 2.303, 2.31, 2.319, 
    2.328, 2.337, 2.347, 2.357, 2.366, 2.374, 2.381, 2.387, 2.39, 2.393, 
    2.394, 2.393, 2.392, 2.391, 2.388, 2.385, 2.382, 2.378, 2.372, 2.364, 
    2.354, 2.34, 2.322, 2.3, 2.274, 2.242, 2.205, 2.164, 2.119, 2.07, 2.019, 
    1.967, 1.913, 1.861, 1.81, 1.76, 1.714, 1.67, 1.63, 1.594, 1.561, 1.533, 
    1.508, 1.486, 1.469, 1.454, 1.443, 1.434, 1.428, 1.424, 1.422, 1.423, 
    1.425, 1.428, 1.432, 1.438, 1.445, 1.452, 1.46, 1.469, 1.477, 1.486, 
    1.496, 1.504, 1.513, 1.521, 1.529, 1.535, 1.54, 1.544, 1.546, 1.547, 
    1.545, 1.542, 1.537, 1.53, 1.521, 1.51, 1.499, 1.486, 1.471, 1.456, 1.44, 
    1.422, 1.404, 1.386, 1.366, 1.346, 1.326, 1.305, 1.284, 1.263, 1.242, 
    1.221, 1.201, 1.181, 1.162, 1.143, 1.125, 1.109, 1.093, 1.078, 1.065, 
    1.052, 1.041, 1.03, 1.021, 1.012, 1.004, 0.997, 0.991, 0.984, 0.979, 
    0.973, 0.968, 0.963, 0.959, 0.954, 0.95, 0.946, 0.942, 0.939, 0.936, 
    0.933, 0.931, 0.929, 0.927, 0.925, 0.924, 0.923, 0.923, 0.922, 0.922, 
    0.922, 0.923, 0.923, 0.924, 0.925, 0.927, 0.928, 0.93, 0.933, 0.935, 
    0.938, 0.941, 0.945, 0.949, 0.953, 0.957, 0.962, 0.967, 0.972, 0.978, 
    0.983, 0.989, 0.995, 1.001, 1.008, 1.014, 1.021, 1.027, 1.034, 1.04, 
    1.047, 1.054, 1.06, 1.067, 1.074, 1.08, 1.087, 1.093, 1.1, 1.106, 1.112, 
    1.119, 1.125, 1.131, 1.137, 1.143, 1.149, 1.154, 1.159, 1.163, 1.168, 
    1.171, 1.175, 1.178, 1.181, 1.184, 1.188, 1.19, 1.194, 1.197, 1.201, 
    1.204, 1.208, 1.212, 1.215, 1.219, 1.223, 1.227, 1.23, 1.234, 1.238, 
    1.242, 1.245, 1.249, 1.253, 1.257, 1.261, 1.265, 1.269, 1.273, 1.277, 
    1.281, 1.285, 1.289, 1.294, 1.298, 1.302, 1.306, 1.311, 1.314, 1.318, 
    1.322, 1.325, 1.329, 1.332, 1.335, 1.338, 1.341, 1.343, 1.345, 1.348, 
    1.35, 1.353, 1.355, 1.357, 1.36, 1.362, 1.364, 1.367, 1.369, 1.371, 
    1.372, 1.373, 1.373, 1.373, 1.372, 1.372, 1.37, 1.369, 1.367, 1.365, 
    1.364, 1.363, 1.363, 1.364, 1.365, 1.366, 1.369, 1.372, 1.376, 1.379, 
    1.383, 1.387, 1.391, 1.394, 1.398, 1.401, 1.405, 1.409, 1.412, 1.415, 
    1.418, 1.422, 1.425, 1.428, 1.431, 1.434, 1.437, 1.439, 1.442, 1.444, 
    1.446, 1.448, 1.45, 1.452, 1.454, 1.456, 1.458, 1.461, 1.463, 1.466, 
    1.469, 1.472, 1.475, 1.478, 1.48, 1.483, 1.485, 1.487, 1.489, 1.491, 
    1.492, 1.492, 1.493, 1.493, 1.493, 1.493, 1.492, 1.492, 1.492, 1.491, 
    1.491, 1.491, 1.492, 1.493, 1.493, 1.495, 1.496, 1.499, 1.501, 1.503, 
    1.506, 1.509, 1.512, 1.515, 1.517, 1.519, 1.519, 1.519, 1.517, 1.514, 
    1.51, 1.505, 1.5, 1.494, 1.489, 1.483, 1.479, 1.476, 1.474, 1.474, 1.474, 
    1.476, 1.479, 1.482, 1.485, 1.488, 1.489, 1.489, 1.488, 1.484, 1.479, 
    1.473, 1.466, 1.458, 1.451, 1.444, 1.438, 1.433, 1.431, 1.43, 1.431, 
    1.434, 1.438, 1.444, 1.451, 1.46, 1.468, 1.477, 1.485, 1.494, 1.502, 
    1.509, 1.515, 1.521, 1.527, 1.531, 1.535, 1.539, 1.543, 1.546, 1.548, 
    1.551, 1.553, 1.555, 1.557, 1.558, 1.56, 1.562, 1.563, 1.565, 1.566, 
    1.568, 1.571, 1.573, 1.576, 1.579, 1.582, 1.586, 1.589, 1.593, 1.597, 
    1.601, 1.605, 1.608, 1.612, 1.616, 1.619, 1.623, 1.626, 1.63, 1.633, 
    1.637, 1.641, 1.644, 1.648, 1.651, 1.655, 1.659, 1.663, 1.666, 1.67, 
    1.674, 1.677, 1.681, 1.684, 1.688, 1.692, 1.695, 1.699, 1.703, 1.706, 
    1.71, 1.714, 1.718, 1.721, 1.725, 1.729, 1.732, 1.736, 1.739, 1.743, 
    1.747, 1.751, 1.756, 1.761, 1.766, 1.771, 1.776, 1.782, 1.788, 1.794, 
    1.799, 1.805, 1.809, 1.814, 1.818, 1.821, 1.823, 1.825, 1.825, 1.826, 
    1.825, 1.824, 1.822, 1.82, 1.818, 1.815, 1.813, 1.811, 1.808, 1.807, 
    1.805, 1.804, 1.803, 1.803, 1.803, 1.803, 1.804, 1.805, 1.807, 1.809, 
    1.811, 1.814, 1.817, 1.82, 1.824, 1.828, 1.833, 1.838, 1.843, 1.849, 
    1.855, 1.862, 1.868, 1.876, 1.883, 1.891, 1.899, 1.908, 1.917, 1.927, 
    1.937, 1.947, 1.958, 1.969, 1.98, 1.991, 2.003, 2.015, 2.027, 2.039, 
    2.052, 2.064, 2.076, 2.089, 2.101, 2.114, 2.126, 2.139, 2.151, 2.163, 
    2.175, 2.187, 2.198, 2.209, 2.22, 2.231, 2.241, 2.25, 2.258, 2.266, 
    2.273, 2.279, 2.284, 2.288, 2.291, 2.292, 2.294, 2.294, 2.293, 2.292, 
    2.29, 2.288, 2.285, 2.281, 2.277, 2.273, 2.268, 2.262, 2.256, 2.249, 
    2.242, 2.233, 2.224, 2.214, 2.204, 2.192, 2.181, 2.168, 2.155, 2.142, 
    2.128, 2.115, 2.101, 2.086, 2.072, 2.057, 2.042, 2.028, 2.012, 1.997, 
    1.981, 1.965, 1.948, 1.931, 1.913, 1.895, 1.876, 1.856, 1.835, 1.812, 
    1.789, 1.764, 1.738, 1.711, 1.683, 1.653, 1.623, 1.592, 1.56, 1.528, 
    1.495, 1.463, 1.431, 1.4, 1.37, 1.34, 1.312, 1.285, 1.26, 1.236, 1.213, 
    1.192, 1.172, 1.154, 1.137, 1.122, 1.108, 1.095, 1.083, 1.072, 1.062, 
    1.053, 1.045, 1.037, 1.03, 1.023, 1.017, 1.011, 1.005, 0.999, 0.993, 
    0.987, 0.982, 0.976, 0.971, 0.965, 0.96, 0.955, 0.95, 0.945, 0.94, 0.935, 
    0.93, 0.924, 0.919, 0.914, 0.908, 0.902, 0.896, 0.889, 0.882, 0.875, 
    0.868, 0.861, 0.853, 0.846, 0.839, 0.831, 0.824, 0.817, 0.81, 0.803, 
    0.797, 0.79, 0.785, 0.779, 0.774, 0.769, 0.764, 0.76, 0.755, 0.751, 
    0.748, 0.744, 0.741, 0.738, 0.735, 0.732, 0.729, 0.727, 0.724, 0.722, 
    0.719, 0.717, 0.715, 0.712, 0.71, 0.708, 0.706, 0.704, 0.702, 0.7, 0.697, 
    0.695, 0.693, 0.691, 0.69, 0.688, 0.686, 0.685, 0.683, 0.682, 0.68, 
    0.679, 0.678, 0.677, 0.677, 0.676, 0.676, 0.677, 0.678, 0.679, 0.681, 
    0.684, 0.688, 0.692, 0.698, 0.703, 0.71, 0.716, 0.723, 0.729, 0.734, 
    0.739, 0.742, 0.745, 0.747, 0.747, 0.747, 0.746, 0.745, 0.744, 0.743, 
    0.742, 0.742, 0.743, 0.744, 0.747, 0.749, 0.752, 0.756, 0.76, 0.764, 
    0.768, 0.772, 0.776, 0.78, 0.784, 0.788, 0.793, 0.797, 0.801, 0.805, 
    0.808, 0.812, 0.816, 0.82, 0.824, 0.827, 0.831, 0.834, 0.837, 0.84, 
    0.843, 0.846, 0.849, 0.852, 0.855, 0.858, 0.861, 0.864, 0.867, 0.871, 
    0.874, 0.878, 0.882, 0.886, 0.889, 0.893, 0.897, 0.9, 0.903, 0.907, 0.91, 
    0.914, 0.917, 0.921, 0.925, 0.928, 0.932, 0.936, 0.94, 0.944, 0.948, 
    0.952, 0.957, 0.96, 0.964, 0.968, 0.971, 0.974, 0.978, 0.981, 0.984, 
    0.987, 0.99, 0.994, 0.997, 1, 1.004, 1.008, 1.01, 1.014, 1.017, 1.02, 
    1.023, 1.025, 1.027, 1.028, 1.03, 1.03, 1.032, 1.033, 1.035, 1.036, 
    1.038, 1.04, 1.042, 1.045, 1.048, 1.051, 1.053, 1.057, 1.06, 1.063, 
    1.066, 1.068, 1.071, 1.072, 1.075, 1.077, 1.079, 1.082, 1.084, 1.086, 
    1.089, 1.091, 1.093, 1.095, 1.097, 1.099, 1.101, 1.101, 1.102, 1.104, 
    1.104, 1.105, 1.106, 1.107, 1.109, 1.11, 1.112, 1.114, 1.116, 1.118, 
    1.12, 1.122, 1.125, 1.126, 1.127, 1.129, 1.13, 1.131, 1.132, 1.133, 
    1.134, 1.135, 1.135, 1.136, 1.138, 1.139, 1.14, 1.141, 1.142, 1.143, 
    1.144, 1.145, 1.146, 1.147, 1.148, 1.15, 1.151, 1.153, 1.154, 1.156, 
    1.157, 1.158, 1.159, 1.16, 1.162, 1.162, 1.163, 1.164, 1.165, 1.165, 
    1.166, 1.167, 1.168, 1.169, 1.171, 1.171, 1.173, 1.174, 1.175, 1.177, 
    1.177, 1.179, 1.179, 1.181, 1.181, 1.183, 1.183, 1.185, 1.185, 1.186, 
    1.187, 1.188, 1.189, 1.19, 1.191, 1.192, 1.193, 1.194, 1.194, 1.195, 
    1.196, 1.197, 1.198, 1.198, 1.199, 1.2, 1.201, 1.201, 1.202, 1.203, 
    1.204, 1.204, 1.205, 1.205, 1.206, 1.207, 1.207, 1.208, 1.208, 1.209, 
    1.209, 1.21, 1.211, 1.211, 1.211, 1.212, 1.212, 1.213, 1.213, 1.214, 
    1.214, 1.215, 1.215, 1.216, 1.217, 1.217, 1.218, 1.218, 1.218, 1.219, 
    1.219, 1.22, 1.22, 1.221, 1.221, 1.221, 1.222, 1.222, 1.222, 1.223, 
    1.223, 1.224, 1.224, 1.225, 1.225, 1.225, 1.226, 1.226, 1.226, 1.226, 
    1.227, 1.227, 1.228, 1.228, 1.228, 1.228, 1.229, 1.229, 1.229, 1.23, 
    1.23, 1.23, 1.231, 1.231, 1.231, 1.231, 1.232, 1.232, 1.233, 1.233, 
    1.233, 1.233, 1.234, 1.234, 1.235, 1.234, 1.235, 1.235, 1.235, 1.235, 
    1.236, 1.236, 1.236, 1.237, 1.237, 1.237, 1.237, 1.237, 1.237, 1.238, 
    1.238, 1.238, 1.239, 1.239, 1.239, 1.24, 1.24, 1.24, 1.24, 1.241, 1.241, 
    1.242, 1.242, 1.242, 1.242, 1.243, 1.243, 1.244, 1.244, 1.244, 1.244, 
    1.244, 1.244, 1.245, 1.245, 1.245, 1.245, 1.246, 1.246, 1.246, 1.247, 
    1.247, 1.247, 1.247, 1.248, 1.248, 1.249, 1.249, 1.249, 1.249, 1.25, 
    1.25, 1.251, 1.251, 1.251, 1.251, 1.251, 1.252, 1.252, 1.253, 1.253, 
    1.253, 1.254, 1.254, 1.255, 1.255, 1.255, 1.255, 1.256, 1.256, 1.256, 
    1.257, 1.257, 1.257, 1.258, 1.258, 1.258, 1.258, 1.258, 1.259, 1.259, 
    1.26, 1.26, 1.26, 1.261, 1.261, 1.262, 1.262, 1.262, 1.263, 1.263, 1.263, 
    1.264, 1.264, 1.265, 1.265, 1.265, 1.266, 1.266, 1.266, 1.266, 1.267, 
    1.267, 1.268, 1.268, 1.268, 1.269, 1.269, 1.269, 1.27, 1.27, 1.27, 1.271, 
    1.271, 1.271, 1.272, 1.272, 1.273, 1.273, 1.273, 1.273, 1.274, 1.274, 
    1.274, 1.275, 1.275, 1.275, 1.276, 1.276, 1.276, 1.277, 1.277, 1.278, 
    1.278, 1.278, 1.278, 1.279, 1.279, 1.279, 1.279, 1.28, 1.28, 1.28, 1.28, 
    1.281, 1.281, 1.281, 1.282, 1.282, 1.282, 1.282, 1.283, 1.283, 1.283, 
    1.284, 1.284, 1.284, 1.285, 1.285, 1.285, 1.285, 1.286, 1.286, 1.286, 
    1.287, 1.287, 1.287, 1.287, 1.288, 1.288, 1.288, 1.288, 1.289, 1.289, 
    1.289, 1.289, 1.289, 1.29, 1.29, 1.29, 1.29, 1.291, 1.291, 1.291, 1.291, 
    1.292, 1.292, 1.292, 1.292, 1.293, 1.293, 1.293, 1.293, 1.293, 1.293, 
    1.293, 1.294, 1.294, 1.294, 1.294, 1.294, 1.294, 1.295, 1.295, 1.295, 
    1.295, 1.295, 1.296, 1.296, 1.296, 1.296, 1.296, 1.297, 1.297, 1.297, 
    1.297, 1.297, 1.297, 1.298, 1.298, 1.298, 1.298, 1.299, 1.299, 1.299, 
    1.299, 1.299, 1.3, 1.3, 1.3, 1.3, 1.3, 1.301, 1.301, 1.301, 1.301, 1.301, 
    1.301, 1.302, 1.302, 1.302, 1.302, 1.302, 1.302, 1.303, 1.303, 1.303, 
    1.303, 1.303, 1.303, 1.304, 1.304, 1.304, 1.304, 1.304, 1.304, 1.304, 
    1.305, 1.305, 1.305, 1.305, 1.305, 1.305, 1.305, 1.305, 1.305, 1.305, 
    1.306, 1.306, 1.306, 1.306, 1.306, 1.307, 1.307, 1.307, 1.307, 1.307, 
    1.308, 1.308, 1.308, 1.308, 1.308, 1.308, 1.309, 1.309, 1.309, 1.309, 
    1.309, 1.309, 1.309, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.311, 1.311, 1.311, 1.311, 1.311, 1.311, 1.312, 1.312, 1.312, 
    1.312, 1.312, 1.312, 1.312, 1.313, 1.313, 1.313, 1.313, 1.313, 1.314, 
    1.314, 1.314, 1.314, 1.314, 1.314, 1.314, 1.315, 1.315, 1.315, 1.315, 
    1.315, 1.315, 1.315, 1.315, 1.316, 1.316, 1.316, 1.316, 1.316, 1.316, 
    1.316, 1.316, 1.317, 1.317, 1.317, 1.317, 1.317, 1.317, 1.317, 1.317, 
    1.318, 1.318, 1.318, 1.318, 1.318, 1.318, 1.319, 1.319, 1.319, 1.319, 
    1.319, 1.319, 1.319, 1.319, 1.319, 1.319, 1.319, 1.319, 1.319, 1.319, 
    1.319, 1.32, 1.32, 1.32, 1.32, 1.32, 1.32, 1.32, 1.32, 1.321, 1.321, 
    1.321, 1.321, 1.321, 1.321, 1.321, 1.321, 1.322, 1.322, 1.322, 1.322, 
    1.322, 1.322, 1.322, 1.322, 1.322, 1.322, 1.322, 1.322, 1.323, 1.323, 
    1.323, 1.323, 1.324, 1.324, 1.324, 1.324, 1.324, 1.324, 1.324, 1.324, 
    1.324, 1.324, 1.324, 1.324, 1.324, 1.325, 1.325, 1.325, 1.325, 1.325, 
    1.325, 1.325, 1.325, 1.325, 1.325, 1.326, 1.326, 1.326, 1.326, 1.326, 
    1.326, 1.326, 1.326, 1.327, 1.327, 1.327, 1.327, 1.327, 1.327, 1.327, 
    1.328, 1.328, 1.328, 1.328, 1.328, 1.328, 1.329, 1.329, 1.329, 1.329, 
    1.329, 1.329, 1.329, 1.329, 1.329, 1.33, 1.33, 1.33, 1.33, 1.33, 1.33, 
    1.33, 1.33, 1.331, 1.331, 1.331, 1.331, 1.331, 1.331, 1.331, 1.332, 
    1.332, 1.332, 1.332, 1.332, 1.332, 1.332, 1.332, 1.333, 1.333, 1.333, 
    1.333, 1.333, 1.333, 1.333, 1.334, 1.334, 1.334, 1.334, 1.334, 1.334, 
    1.334, 1.334, 1.334, 1.334, 1.335, 1.335, 1.335, 1.335, 1.335, 1.335, 
    1.336, 1.336, 1.336, 1.336, 1.336, 1.336, 1.336, 1.337, 1.337, 1.337, 
    1.337, 1.337, 1.338, 1.338, 1.338, 1.338, 1.338, 1.338, 1.339, 1.339, 
    1.339, 1.339, 1.339, 1.339, 1.339, 1.34, 1.339, 1.339, 1.34, 1.34, 1.34, 
    1.34, 1.34, 1.34, 1.34, 1.34, 1.341, 1.341, 1.341, 1.341, 1.341, 1.341, 
    1.341, 1.341, 1.342, 1.342, 1.342, 1.342, 1.342, 1.343, 1.343, 1.343, 
    1.343, 1.343, 1.343, 1.344, 1.344, 1.344, 1.344, 1.344, 1.344, 1.344, 
    1.344, 1.344, 1.345, 1.345, 1.345, 1.345, 1.345, 1.345, 1.346, 1.346, 
    1.346, 1.346, 1.346, 1.346, 1.346, 1.347, 1.347, 1.347, 1.347, 1.347, 
    1.347, 1.348, 1.348, 1.348, 1.348, 1.348, 1.348, 1.348, 1.348, 1.348, 
    1.349, 1.349, 1.349, 1.349, 1.349, 1.35, 1.35, 1.35, 1.35, 1.35, 1.35, 
    1.35, 1.351, 1.351, 1.351, 1.351, 1.351, 1.351, 1.351, 1.351, 1.352, 
    1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 1.352, 1.353, 
    1.353, 1.353, 1.353, 1.353, 1.353, 1.353, 1.354, 1.354, 1.354, 1.354, 
    1.354, 1.354, 1.354, 1.354, 1.354, 1.354, 1.355, 1.355, 1.355, 1.355, 
    1.355, 1.355, 1.355, 1.355, 1.355, 1.355, 1.356, 1.355, 1.355, 1.355, 
    1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 1.356, 
    1.356, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 1.357, 
    1.357, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 1.358, 
    1.358, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 
    1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 1.359, 
    1.359, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 1.36, 
    1.36, 1.36, 1.36, 1.36, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 
    1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 1.361, 
    1.361, 1.361, 1.361, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 
    1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 1.362, 
    1.362, 1.362, 1.362, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 
    1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 1.363, 
    1.363, 1.363, 1.363, 1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 
    1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 1.364, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.372, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 1.375, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 1.374, 
    1.374, 1.374, 1.374, 1.374, 1.374, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 1.372, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 1.371, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 
    1.37, 1.37, 1.37, 1.37, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.366, 1.366, 
    1.366, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 
    1.365, 1.365, 1.365, 1.365, 1.365, 1.365, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 1.366, 
    1.366, 1.366, 1.366, 1.366, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.367, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 
    1.368, 1.368, 1.368, 1.368, 1.369, 1.369, 1.369, 1.369, 1.369, 1.369, 
    1.369, 1.369, 1.369, 1.369, 1.369, 1.37, 1.37, 1.37, 1.37, 1.37, 1.369, 
    1.369, 1.368, 1.368, 1.368, 1.367, 1.367, 1.367, 1.367, 1.367, 1.368, 
    1.368, 1.369, 1.37, 1.37, 1.37, 1.371, 1.371, 1.371, 1.371, 1.371, 1.37, 
    1.37, 1.369, 1.369, 1.369, 1.368, 1.368, 1.368, 1.368, 1.368, 1.369, 
    1.369, 1.37, 1.371, 1.371, 1.372, 1.372, 1.373, 1.373, 1.373, 1.374, 
    1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.373, 1.372, 1.372, 1.371, 
    1.371, 1.371, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.37, 1.371, 1.371, 
    1.372, 1.372, 1.373, 1.373, 1.374, 1.374, 1.374, 1.375, 1.375, 1.375, 
    1.376, 1.376, 1.376, 1.377, 1.377, 1.378, 1.378, 1.378, 1.378, 1.379, 
    1.378, 1.378, 1.378, 1.378, 1.377, 1.376, 1.376, 1.375, 1.374, 1.373, 
    1.372, 1.371, 1.371, 1.37, 1.369, 1.369, 1.368, 1.368, 1.368, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.366, 1.365, 1.365, 1.364, 1.362, 1.361, 
    1.36, 1.358, 1.357, 1.356, 1.355, 1.354, 1.353, 1.353, 1.353, 1.352, 
    1.352, 1.352, 1.351, 1.35, 1.349, 1.348, 1.347, 1.345, 1.344, 1.343, 
    1.342, 1.34, 1.34, 1.339, 1.339, 1.338, 1.338, 1.339, 1.339, 1.34, 1.34, 
    1.341, 1.342, 1.342, 1.343, 1.343, 1.343, 1.343, 1.342, 1.342, 1.341, 
    1.34, 1.34, 1.339, 1.338, 1.338, 1.338, 1.338, 1.339, 1.339, 1.34, 1.341, 
    1.342, 1.343, 1.344, 1.345, 1.345, 1.346, 1.346, 1.346, 1.346, 1.346, 
    1.346, 1.346, 1.346, 1.346, 1.347, 1.348, 1.349, 1.349, 1.35, 1.352, 
    1.353, 1.353, 1.354, 1.354, 1.355, 1.355, 1.355, 1.355, 1.356, 1.356, 
    1.356, 1.357, 1.357, 1.358, 1.358, 1.358, 1.359, 1.36, 1.36, 1.361, 
    1.362, 1.363, 1.363, 1.364, 1.365, 1.365, 1.366, 1.366, 1.367, 1.367, 
    1.367, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.368, 1.367, 
    1.367, 1.367, 1.367, 1.367, 1.368, 1.368, 1.369, 1.369, 1.37, 1.371, 
    1.372, 1.373, 1.374, 1.375, 1.376, 1.377, 1.378, 1.378, 1.379, 1.379, 
    1.379, 1.38, 1.38, 1.379, 1.379, 1.378, 1.378, 1.378, 1.377, 1.377, 
    1.377, 1.377, 1.377, 1.377, 1.377, 1.377, 1.378, 1.378, 1.378, 1.378, 
    1.379, 1.379, 1.379, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 1.378, 
    1.378, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.379, 1.378, 1.378, 
    1.378, 1.378, 1.377, 1.377, 1.377, 1.377, 1.378, 1.378, 1.379, 1.379, 
    1.38, 1.381, 1.381, 1.382, 1.382, 1.382, 1.382, 1.381, 1.381, 1.38, 
    1.379, 1.378, 1.378, 1.378, 1.378, 1.378, 1.379, 1.38, 1.382, 1.382, 
    1.383, 1.384, 1.384, 1.384, 1.383, 1.382, 1.381, 1.379, 1.378, 1.377, 
    1.376, 1.375, 1.375, 1.375, 1.376, 1.377, 1.378, 1.379, 1.38, 1.381, 
    1.382, 1.382, 1.382, 1.382, 1.382, 1.382, 1.381, 1.381, 1.381, 1.381, 
    1.382, 1.382, 1.382, 1.383, 1.383, 1.383, 1.383, 1.383, 1.382, 1.382, 
    1.381, 1.381, 1.38, 1.38, 1.38, 1.38, 1.381, 1.382, 1.382, 1.383, 1.383, 
    1.384, 1.384, 1.384, 1.384, 1.383, 1.383, 1.382, 1.381, 1.381, 1.381, 
    1.381, 1.38, 1.38, 1.381, 1.381, 1.381, 1.381, 1.381, 1.381, 1.381, 
    1.381, 1.381, 1.38, 1.38, 1.38, 1.38, 1.38, 1.38, 1.381, 1.382, 1.382, 
    1.383, 1.384, 1.384, 1.385, 1.385, 1.385, 1.384, 1.384, 1.383, 1.382, 
    1.382, 1.381, 1.381, 1.381, 1.381, 1.381, 1.381, 1.381, 1.382, 1.382, 
    1.382, 1.382, 1.383, 1.383, 1.384, 1.384, 1.385, 1.385, 1.385, 1.385, 
    1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 
    1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.385, 1.384, 1.384, 
    1.384, 1.384, 1.384, 1.384, 1.384, 1.383, 1.383, 1.382, 1.382, 1.381, 
    1.381, 1.38, 1.38, 1.38, 1.38, 1.38, 1.38, 1.38, 1.38, 1.38, 1.38, 1.381, 
    1.381, 1.381, 1.382, 1.382, 1.382, 1.382, 1.382, 1.382, 1.382, 1.381, 
    1.381, 1.381, 1.381, 1.381, 1.381, 1.381, 1.38, 1.38, 1.38, 1.381, 1.381, 
    1.381, 1.381, 1.381, 1.381 ;

 idx_rfr_illite_img = 0.066, 0.064, 0.063, 0.062, 0.061, 0.06, 0.059, 0.059, 
    0.059, 0.06, 0.061, 0.062, 0.062, 0.062, 0.062, 0.063, 0.064, 0.065, 
    0.068, 0.071, 0.075, 0.08, 0.086, 0.091, 0.097, 0.104, 0.113, 0.124, 
    0.136, 0.15, 0.166, 0.183, 0.201, 0.219, 0.235, 0.252, 0.267, 0.282, 
    0.297, 0.311, 0.325, 0.337, 0.349, 0.36, 0.37, 0.379, 0.386, 0.392, 
    0.398, 0.404, 0.409, 0.413, 0.416, 0.419, 0.421, 0.423, 0.423, 0.42, 
    0.415, 0.406, 0.395, 0.382, 0.368, 0.354, 0.34, 0.328, 0.318, 0.311, 
    0.305, 0.3, 0.296, 0.293, 0.29, 0.287, 0.284, 0.283, 0.281, 0.281, 0.28, 
    0.279, 0.278, 0.276, 0.274, 0.271, 0.266, 0.261, 0.255, 0.25, 0.244, 
    0.239, 0.234, 0.23, 0.227, 0.223, 0.22, 0.218, 0.215, 0.212, 0.21, 0.208, 
    0.206, 0.204, 0.202, 0.201, 0.201, 0.2, 0.2, 0.199, 0.198, 0.198, 0.196, 
    0.194, 0.191, 0.188, 0.185, 0.182, 0.18, 0.178, 0.176, 0.175, 0.175, 
    0.176, 0.177, 0.179, 0.181, 0.184, 0.186, 0.189, 0.193, 0.197, 0.201, 
    0.205, 0.209, 0.213, 0.216, 0.218, 0.219, 0.219, 0.218, 0.216, 0.214, 
    0.211, 0.208, 0.205, 0.202, 0.199, 0.196, 0.192, 0.188, 0.184, 0.18, 
    0.176, 0.172, 0.17, 0.167, 0.165, 0.163, 0.162, 0.162, 0.162, 0.162, 
    0.163, 0.164, 0.164, 0.165, 0.165, 0.164, 0.163, 0.162, 0.162, 0.162, 
    0.163, 0.164, 0.165, 0.166, 0.167, 0.167, 0.167, 0.167, 0.168, 0.169, 
    0.171, 0.173, 0.175, 0.177, 0.178, 0.18, 0.183, 0.185, 0.188, 0.191, 
    0.196, 0.201, 0.207, 0.214, 0.221, 0.228, 0.235, 0.242, 0.249, 0.256, 
    0.262, 0.268, 0.274, 0.279, 0.284, 0.288, 0.292, 0.295, 0.297, 0.298, 
    0.298, 0.297, 0.295, 0.292, 0.288, 0.283, 0.277, 0.27, 0.263, 0.256, 
    0.249, 0.242, 0.236, 0.23, 0.225, 0.221, 0.217, 0.214, 0.212, 0.21, 
    0.209, 0.208, 0.207, 0.206, 0.206, 0.206, 0.205, 0.205, 0.205, 0.205, 
    0.205, 0.205, 0.205, 0.206, 0.206, 0.206, 0.207, 0.208, 0.209, 0.21, 
    0.212, 0.213, 0.215, 0.218, 0.22, 0.222, 0.225, 0.228, 0.23, 0.233, 
    0.236, 0.239, 0.241, 0.244, 0.247, 0.25, 0.253, 0.256, 0.258, 0.261, 
    0.263, 0.265, 0.268, 0.27, 0.272, 0.274, 0.277, 0.279, 0.282, 0.284, 
    0.287, 0.29, 0.293, 0.296, 0.299, 0.303, 0.307, 0.312, 0.318, 0.324, 
    0.332, 0.34, 0.349, 0.359, 0.369, 0.379, 0.39, 0.4, 0.41, 0.419, 0.428, 
    0.436, 0.443, 0.449, 0.455, 0.459, 0.464, 0.468, 0.472, 0.477, 0.482, 
    0.488, 0.494, 0.501, 0.508, 0.514, 0.52, 0.525, 0.528, 0.529, 0.528, 
    0.524, 0.518, 0.51, 0.5, 0.488, 0.476, 0.463, 0.451, 0.44, 0.43, 0.422, 
    0.416, 0.414, 0.416, 0.421, 0.429, 0.441, 0.456, 0.472, 0.489, 0.506, 
    0.521, 0.534, 0.543, 0.548, 0.549, 0.546, 0.54, 0.533, 0.524, 0.515, 
    0.507, 0.501, 0.498, 0.499, 0.502, 0.51, 0.521, 0.535, 0.551, 0.57, 0.59, 
    0.61, 0.631, 0.652, 0.672, 0.691, 0.71, 0.729, 0.746, 0.762, 0.777, 
    0.791, 0.804, 0.814, 0.823, 0.83, 0.836, 0.84, 0.843, 0.844, 0.844, 
    0.844, 0.843, 0.842, 0.842, 0.842, 0.843, 0.846, 0.851, 0.857, 0.866, 
    0.877, 0.89, 0.906, 0.923, 0.942, 0.963, 0.984, 1.01, 1.03, 1.05, 1.08, 
    1.1, 1.12, 1.15, 1.18, 1.2, 1.23, 1.27, 1.3, 1.34, 1.37, 1.41, 1.45, 
    1.48, 1.52, 1.55, 1.57, 1.59, 1.61, 1.62, 1.63, 1.62, 1.62, 1.61, 1.59, 
    1.57, 1.55, 1.52, 1.5, 1.47, 1.44, 1.41, 1.38, 1.35, 1.32, 1.29, 1.26, 
    1.24, 1.21, 1.19, 1.17, 1.15, 1.13, 1.12, 1.1, 1.09, 1.08, 1.07, 1.06, 
    1.06, 1.05, 1.05, 1.05, 1.05, 1.06, 1.06, 1.07, 1.08, 1.09, 1.1, 1.11, 
    1.12, 1.13, 1.14, 1.15, 1.17, 1.18, 1.18, 1.19, 1.2, 1.21, 1.21, 1.22, 
    1.22, 1.23, 1.23, 1.23, 1.23, 1.22, 1.22, 1.21, 1.21, 1.2, 1.19, 1.18, 
    1.17, 1.15, 1.14, 1.12, 1.11, 1.1, 1.08, 1.06, 1.05, 1.03, 1.02, 1, 
    0.984, 0.969, 0.954, 0.94, 0.925, 0.911, 0.897, 0.883, 0.869, 0.856, 
    0.842, 0.828, 0.814, 0.8, 0.787, 0.773, 0.759, 0.746, 0.732, 0.719, 
    0.705, 0.692, 0.679, 0.666, 0.653, 0.64, 0.628, 0.615, 0.602, 0.59, 
    0.577, 0.565, 0.552, 0.54, 0.528, 0.516, 0.505, 0.493, 0.482, 0.471, 
    0.46, 0.449, 0.439, 0.429, 0.419, 0.41, 0.401, 0.392, 0.384, 0.376, 
    0.368, 0.361, 0.354, 0.347, 0.341, 0.335, 0.329, 0.324, 0.318, 0.313, 
    0.309, 0.304, 0.3, 0.296, 0.292, 0.288, 0.285, 0.282, 0.28, 0.278, 0.276, 
    0.274, 0.273, 0.271, 0.27, 0.269, 0.267, 0.265, 0.263, 0.261, 0.258, 
    0.256, 0.253, 0.25, 0.248, 0.245, 0.242, 0.24, 0.237, 0.235, 0.233, 0.23, 
    0.228, 0.226, 0.224, 0.221, 0.219, 0.217, 0.215, 0.213, 0.211, 0.21, 
    0.208, 0.206, 0.205, 0.203, 0.202, 0.201, 0.2, 0.199, 0.198, 0.198, 
    0.198, 0.197, 0.198, 0.198, 0.198, 0.198, 0.199, 0.199, 0.2, 0.201, 
    0.201, 0.201, 0.202, 0.202, 0.202, 0.203, 0.203, 0.203, 0.204, 0.205, 
    0.206, 0.207, 0.208, 0.21, 0.212, 0.213, 0.215, 0.216, 0.216, 0.216, 
    0.216, 0.215, 0.213, 0.21, 0.207, 0.203, 0.2, 0.196, 0.192, 0.188, 0.184, 
    0.181, 0.179, 0.176, 0.175, 0.173, 0.172, 0.171, 0.17, 0.169, 0.169, 
    0.169, 0.169, 0.168, 0.168, 0.168, 0.169, 0.169, 0.17, 0.17, 0.171, 
    0.172, 0.172, 0.173, 0.174, 0.174, 0.174, 0.174, 0.174, 0.174, 0.174, 
    0.174, 0.175, 0.175, 0.176, 0.177, 0.178, 0.18, 0.182, 0.184, 0.186, 
    0.188, 0.191, 0.193, 0.195, 0.197, 0.199, 0.201, 0.202, 0.203, 0.204, 
    0.205, 0.205, 0.205, 0.204, 0.204, 0.204, 0.203, 0.202, 0.202, 0.201, 
    0.202, 0.202, 0.203, 0.204, 0.207, 0.21, 0.213, 0.218, 0.223, 0.228, 
    0.233, 0.237, 0.241, 0.244, 0.246, 0.246, 0.245, 0.243, 0.239, 0.235, 
    0.23, 0.225, 0.221, 0.218, 0.215, 0.214, 0.214, 0.216, 0.218, 0.222, 
    0.226, 0.229, 0.231, 0.233, 0.232, 0.23, 0.225, 0.219, 0.211, 0.201, 
    0.191, 0.18, 0.169, 0.158, 0.148, 0.139, 0.131, 0.124, 0.119, 0.115, 
    0.112, 0.111, 0.111, 0.111, 0.112, 0.113, 0.114, 0.116, 0.117, 0.119, 
    0.12, 0.121, 0.123, 0.124, 0.125, 0.126, 0.126, 0.127, 0.127, 0.127, 
    0.126, 0.126, 0.125, 0.124, 0.122, 0.121, 0.12, 0.118, 0.117, 0.116, 
    0.115, 0.114, 0.113, 0.113, 0.113, 0.113, 0.113, 0.113, 0.113, 0.114, 
    0.114, 0.114, 0.114, 0.115, 0.115, 0.115, 0.116, 0.116, 0.117, 0.118, 
    0.119, 0.119, 0.12, 0.121, 0.122, 0.123, 0.124, 0.125, 0.126, 0.127, 
    0.128, 0.129, 0.13, 0.132, 0.133, 0.135, 0.136, 0.137, 0.139, 0.14, 
    0.142, 0.143, 0.144, 0.145, 0.147, 0.148, 0.149, 0.151, 0.153, 0.155, 
    0.158, 0.161, 0.165, 0.17, 0.175, 0.181, 0.187, 0.193, 0.2, 0.207, 0.214, 
    0.22, 0.227, 0.233, 0.239, 0.244, 0.248, 0.252, 0.255, 0.257, 0.259, 
    0.26, 0.26, 0.26, 0.259, 0.259, 0.257, 0.256, 0.255, 0.253, 0.251, 0.249, 
    0.248, 0.246, 0.244, 0.241, 0.239, 0.237, 0.235, 0.233, 0.231, 0.229, 
    0.228, 0.226, 0.225, 0.224, 0.222, 0.222, 0.221, 0.221, 0.22, 0.221, 
    0.221, 0.222, 0.223, 0.225, 0.227, 0.23, 0.233, 0.237, 0.241, 0.246, 
    0.252, 0.258, 0.265, 0.272, 0.28, 0.289, 0.298, 0.308, 0.319, 0.331, 
    0.343, 0.356, 0.369, 0.384, 0.399, 0.415, 0.432, 0.449, 0.468, 0.487, 
    0.507, 0.527, 0.548, 0.569, 0.591, 0.613, 0.635, 0.657, 0.679, 0.7, 
    0.722, 0.743, 0.764, 0.785, 0.807, 0.827, 0.848, 0.869, 0.891, 0.912, 
    0.933, 0.954, 0.974, 0.995, 1.02, 1.04, 1.05, 1.07, 1.09, 1.11, 1.13, 
    1.15, 1.16, 1.18, 1.2, 1.21, 1.23, 1.24, 1.26, 1.27, 1.29, 1.3, 1.32, 
    1.33, 1.35, 1.36, 1.38, 1.39, 1.41, 1.42, 1.44, 1.45, 1.47, 1.48, 1.49, 
    1.5, 1.51, 1.52, 1.53, 1.53, 1.53, 1.53, 1.53, 1.53, 1.52, 1.51, 1.5, 
    1.49, 1.48, 1.47, 1.46, 1.44, 1.42, 1.41, 1.39, 1.38, 1.36, 1.34, 1.33, 
    1.31, 1.3, 1.28, 1.27, 1.25, 1.24, 1.23, 1.21, 1.2, 1.19, 1.18, 1.17, 
    1.16, 1.15, 1.14, 1.13, 1.12, 1.12, 1.11, 1.1, 1.09, 1.09, 1.08, 1.07, 
    1.06, 1.06, 1.05, 1.04, 1.04, 1.03, 1.03, 1.02, 1.02, 1.01, 1, 0.997, 
    0.99, 0.983, 0.975, 0.968, 0.959, 0.951, 0.942, 0.934, 0.924, 0.915, 
    0.906, 0.896, 0.886, 0.877, 0.867, 0.857, 0.848, 0.838, 0.829, 0.819, 
    0.81, 0.8, 0.791, 0.782, 0.773, 0.764, 0.756, 0.747, 0.738, 0.73, 0.721, 
    0.713, 0.704, 0.696, 0.688, 0.679, 0.671, 0.663, 0.654, 0.646, 0.637, 
    0.628, 0.62, 0.611, 0.602, 0.593, 0.584, 0.575, 0.565, 0.556, 0.546, 
    0.537, 0.527, 0.516, 0.506, 0.495, 0.484, 0.473, 0.462, 0.452, 0.441, 
    0.431, 0.421, 0.412, 0.404, 0.398, 0.392, 0.388, 0.384, 0.381, 0.379, 
    0.377, 0.375, 0.373, 0.37, 0.366, 0.361, 0.356, 0.35, 0.343, 0.335, 
    0.327, 0.319, 0.311, 0.303, 0.296, 0.289, 0.282, 0.275, 0.269, 0.264, 
    0.258, 0.253, 0.248, 0.243, 0.238, 0.234, 0.229, 0.225, 0.221, 0.217, 
    0.214, 0.21, 0.206, 0.203, 0.2, 0.197, 0.194, 0.19, 0.187, 0.184, 0.18, 
    0.177, 0.173, 0.17, 0.166, 0.162, 0.159, 0.155, 0.152, 0.148, 0.145, 
    0.142, 0.139, 0.137, 0.134, 0.132, 0.129, 0.126, 0.123, 0.121, 0.118, 
    0.116, 0.113, 0.111, 0.108, 0.106, 0.104, 0.102, 0.1, 0.098, 0.097, 
    0.096, 0.094, 0.094, 0.093, 0.092, 0.091, 0.09, 0.088, 0.088, 0.086, 
    0.086, 0.085, 0.084, 0.083, 0.083, 0.082, 0.082, 0.083, 0.082, 0.083, 
    0.084, 0.084, 0.084, 0.085, 0.083, 0.083, 0.082, 0.081, 0.08, 0.078, 
    0.076, 0.074, 0.073, 0.071, 0.071, 0.069, 0.068, 0.068, 0.068, 0.068, 
    0.068, 0.068, 0.068, 0.067, 0.068, 0.067, 0.067, 0.068, 0.067, 0.067, 
    0.067, 0.068, 0.068, 0.069, 0.069, 0.071, 0.071, 0.071, 0.071, 0.072, 
    0.071, 0.071, 0.07, 0.069, 0.068, 0.067, 0.067, 0.066, 0.066, 0.066, 
    0.066, 0.067, 0.068, 0.068, 0.069, 0.069, 0.07, 0.07, 0.07, 0.07, 0.07, 
    0.07, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.068, 0.068, 
    0.068, 0.067, 0.067, 0.067, 0.066, 0.066, 0.066, 0.066, 0.067, 0.067, 
    0.067, 0.067, 0.067, 0.068, 0.068, 0.068, 0.067, 0.067, 0.067, 0.067, 
    0.067, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 0.066, 
    0.066, 0.066, 0.066, 0.066, 0.066, 0.067, 0.067, 0.067, 0.067, 0.067, 
    0.067, 0.067, 0.067, 0.068, 0.068, 0.068, 0.068, 0.068, 0.068, 0.069, 
    0.069, 0.069, 0.069, 0.069, 0.07, 0.07, 0.07, 0.07, 0.07, 0.071, 0.071, 
    0.071, 0.071, 0.071, 0.071, 0.071, 0.072, 0.072, 0.072, 0.072, 0.072, 
    0.072, 0.072, 0.072, 0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 0.073, 
    0.073, 0.073, 0.073, 0.073, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 
    0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 
    0.074, 0.074, 0.074, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.074, 0.075, 0.074, 0.074, 
    0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 
    0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.074, 0.073, 0.074, 0.073, 
    0.073, 0.073, 0.073, 0.073, 0.072, 0.072, 0.072, 0.072, 0.072, 0.072, 
    0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.071, 0.07, 0.07, 0.07, 0.07, 
    0.07, 0.07, 0.07, 0.07, 0.07, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 
    0.069, 0.068, 0.068, 0.068, 0.067, 0.067, 0.067, 0.067, 0.067, 0.067, 
    0.066, 0.066, 0.066, 0.066, 0.066, 0.065, 0.065, 0.065, 0.065, 0.065, 
    0.065, 0.064, 0.064, 0.064, 0.064, 0.064, 0.063, 0.063, 0.063, 0.063, 
    0.063, 0.063, 0.063, 0.063, 0.062, 0.062, 0.062, 0.062, 0.062, 0.062, 
    0.062, 0.061, 0.061, 0.061, 0.061, 0.06, 0.06, 0.06, 0.06, 0.06, 0.06, 
    0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.058, 
    0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 0.057, 0.057, 
    0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.057, 0.056, 
    0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 0.056, 
    0.055, 0.056, 0.056, 0.056, 0.056, 0.055, 0.056, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 0.055, 
    0.055, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.055, 0.055, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 
    0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.054, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 
    0.052, 0.053, 0.053, 0.052, 0.053, 0.053, 0.053, 0.053, 0.052, 0.052, 
    0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.052, 0.051, 0.052, 0.052, 
    0.051, 0.052, 0.052, 0.051, 0.051, 0.052, 0.051, 0.051, 0.052, 0.051, 
    0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 
    0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 0.051, 
    0.051, 0.051, 0.051, 0.051, 0.051, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.049, 0.05, 0.05, 0.05, 0.049, 0.049, 0.05, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.048, 0.048, 0.049, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.047, 0.048, 0.048, 0.048, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.045, 0.045, 
    0.046, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.043, 0.043, 0.044, 0.044, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.04, 0.041, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.039, 0.039, 0.04, 0.04, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.038, 0.038, 0.038, 0.038, 0.039, 0.038, 0.038, 0.039, 
    0.038, 0.038, 0.039, 0.039, 0.038, 0.039, 0.039, 0.039, 0.039, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.039, 0.039, 0.039, 0.038, 0.038, 0.038, 0.038, 0.038, 0.039, 
    0.038, 0.038, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.04, 0.04, 0.04, 0.039, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.041, 0.041, 0.04, 0.04, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.042, 0.042, 0.042, 0.041, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.042, 0.042, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.042, 0.042, 0.043, 
    0.043, 0.043, 0.042, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.044, 0.044, 0.044, 0.044, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.043, 0.043, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.043, 0.043, 0.044, 
    0.044, 0.044, 0.043, 0.043, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.043, 0.043, 0.044, 0.044, 0.044, 0.043, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.044, 0.044, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.045, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.046, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.048, 0.048, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.047, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.05, 0.05, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.049, 0.049, 0.049, 0.05, 0.05, 0.05, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 0.049, 
    0.049, 0.049, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.049, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 0.046, 
    0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.045, 0.045, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.045, 0.045, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.044, 
    0.044, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.042, 0.042, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.04, 0.04, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.039, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.037, 0.037, 0.037, 0.037, 
    0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 
    0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.036, 0.036, 0.036, 
    0.036, 0.037, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 
    0.036, 0.036, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 
    0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.034, 0.034, 0.034, 
    0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 
    0.034, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 
    0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.033, 0.032, 0.032, 
    0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 0.032, 
    0.032, 0.032, 0.032, 0.032, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.029, 0.029, 0.029, 0.029, 0.029, 
    0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 0.029, 
    0.029, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 
    0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 
    0.028, 0.028, 0.028, 0.028, 0.028, 0.028, 0.027, 0.027, 0.027, 0.027, 
    0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 
    0.027, 0.027, 0.027, 0.026, 0.026, 0.027, 0.026, 0.026, 0.026, 0.026, 
    0.026, 0.026, 0.026, 0.027, 0.027, 0.027, 0.027, 0.027, 0.028, 0.028, 
    0.028, 0.028, 0.028, 0.028, 0.028, 0.027, 0.027, 0.026, 0.026, 0.025, 
    0.025, 0.025, 0.024, 0.024, 0.025, 0.025, 0.025, 0.026, 0.027, 0.027, 
    0.027, 0.028, 0.028, 0.028, 0.028, 0.027, 0.027, 0.026, 0.026, 0.025, 
    0.025, 0.024, 0.024, 0.023, 0.023, 0.023, 0.024, 0.024, 0.024, 0.025, 
    0.025, 0.026, 0.026, 0.027, 0.027, 0.027, 0.028, 0.028, 0.029, 0.029, 
    0.029, 0.029, 0.029, 0.029, 0.029, 0.028, 0.028, 0.027, 0.027, 0.026, 
    0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 
    0.027, 0.027, 0.027, 0.027, 0.028, 0.028, 0.028, 0.029, 0.03, 0.03, 
    0.031, 0.032, 0.033, 0.034, 0.035, 0.036, 0.037, 0.038, 0.039, 0.039, 
    0.04, 0.04, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.042, 0.042, 0.043, 0.043, 0.044, 0.044, 
    0.045, 0.046, 0.046, 0.046, 0.046, 0.045, 0.045, 0.044, 0.043, 0.043, 
    0.042, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.04, 0.039, 0.038, 0.037, 0.036, 0.034, 0.033, 0.031, 0.03, 0.028, 
    0.027, 0.025, 0.024, 0.023, 0.022, 0.022, 0.022, 0.021, 0.021, 0.022, 
    0.022, 0.022, 0.021, 0.021, 0.021, 0.02, 0.019, 0.017, 0.016, 0.014, 
    0.013, 0.011, 0.01, 0.009, 0.008, 0.007, 0.006, 0.006, 0.006, 0.006, 
    0.006, 0.006, 0.006, 0.005, 0.005, 0.004, 0.003, 0.002, 0.001, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001, 0.001, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.002, 0.002, 0.002, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.005, 0.005, 0.005, 0.005, 0.005, 0.004, 0.004, 0.003, 
    0.003, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.003, 0.003, 0.004, 
    0.005, 0.005, 0.006, 0.006, 0.006, 0.007, 0.006, 0.005, 0.005, 0.004, 
    0.003, 0.003, 0.002, 0.002, 0.003, 0.004, 0.005, 0.006, 0.007, 0.009, 
    0.01, 0.01, 0.01, 0.01, 0.009, 0.008, 0.007, 0.006, 0.004, 0.003, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.003, 0.004, 0.004, 0.005, 0.005, 
    0.005, 0.005, 0.005, 0.004, 0.004, 0.004, 0.004, 0.005, 0.005, 0.006, 
    0.006, 0.007, 0.007, 0.007, 0.007, 0.007, 0.006, 0.006, 0.006, 0.005, 
    0.004, 0.004, 0.004, 0.004, 0.005, 0.005, 0.006, 0.006, 0.007, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.007, 0.007, 0.006, 0.006, 0.006, 
    0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.005, 
    0.005, 0.004, 0.004, 0.003, 0.003, 0.003, 0.003, 0.004, 0.004, 0.005, 
    0.005, 0.006, 0.007, 0.007, 0.008, 0.008, 0.007, 0.007, 0.007, 0.006, 
    0.006, 0.005, 0.005, 0.004, 0.004, 0.004, 0.004, 0.003, 0.003, 0.003, 
    0.003, 0.003, 0.004, 0.004, 0.004, 0.005, 0.005, 0.005, 0.006, 0.006, 
    0.006, 0.006, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 
    0.007, 0.008, 0.008, 0.008, 0.008, 0.008, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.01, 0.01, 0.01, 0.01, 0.01, 0.009, 0.009, 0.008, 0.008, 0.008, 
    0.007, 0.007, 0.007, 0.006, 0.006, 0.006, 0.005, 0.005, 0.005, 0.005, 
    0.005, 0.005, 0.005, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 
    0.006, 0.006, 0.006, 0.005, 0.005, 0.005, 0.004, 0.005, 0.004, 0.004, 
    0.004, 0.004 ;

 idx_rfr_illite_rl_ee = 0.02, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.011, 
    0.011, 0.011, 0.012, 0.012, 0.012, 0.013, 0.013, 0.014, 0.015, 0.016, 
    0.016, 0.017, 0.018, 0.019, 0.02, 0.021, 0.021, 0.022, 0.023, 0.023, 
    0.024, 0.024, 0.025, 0.025, 0.025, 0.025, 0.026, 0.026, 0.026, 0.026, 
    0.026, 0.026, 0.026, 0.026, 0.026, 0.025, 0.025, 0.025, 0.024, 0.024, 
    0.023, 0.022, 0.022, 0.021, 0.021, 0.02, 0.02, 0.02, 0.019, 0.019, 0.019, 
    0.019, 0.019, 0.019, 0.019, 0.019, 0.019, 0.019, 0.019, 0.018, 0.018, 
    0.018, 0.018, 0.018, 0.018, 0.017, 0.017, 0.017, 0.017, 0.017, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.016, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 
    0.016, 0.016, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.014, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.016, 0.016, 
    0.016, 0.016, 0.017, 0.017, 0.017, 0.018, 0.018, 0.018, 0.019, 0.019, 
    0.019, 0.019, 0.019, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 
    0.02, 0.019, 0.019, 0.019, 0.019, 0.018, 0.018, 0.018, 0.018, 0.017, 
    0.017, 0.017, 0.017, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.017, 0.017, 0.017, 
    0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.018, 0.018, 0.018, 0.018, 
    0.018, 0.018, 0.019, 0.019, 0.019, 0.019, 0.019, 0.019, 0.019, 0.019, 
    0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.021, 0.021, 0.021, 0.021, 
    0.021, 0.021, 0.022, 0.022, 0.022, 0.022, 0.023, 0.023, 0.024, 0.024, 
    0.025, 0.025, 0.026, 0.026, 0.027, 0.027, 0.027, 0.028, 0.028, 0.028, 
    0.029, 0.029, 0.029, 0.029, 0.029, 0.03, 0.03, 0.03, 0.03, 0.03, 0.031, 
    0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.031, 0.03, 0.03, 
    0.029, 0.029, 0.028, 0.028, 0.027, 0.027, 0.027, 0.026, 0.026, 0.026, 
    0.027, 0.027, 0.028, 0.028, 0.029, 0.03, 0.031, 0.032, 0.032, 0.033, 
    0.033, 0.033, 0.033, 0.033, 0.033, 0.032, 0.032, 0.031, 0.031, 0.031, 
    0.031, 0.031, 0.032, 0.032, 0.033, 0.034, 0.035, 0.036, 0.037, 0.038, 
    0.04, 0.041, 0.042, 0.043, 0.043, 0.044, 0.045, 0.046, 0.046, 0.047, 
    0.047, 0.047, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.047, 
    0.047, 0.047, 0.047, 0.047, 0.048, 0.048, 0.048, 0.049, 0.049, 0.05, 
    0.051, 0.052, 0.053, 0.054, 0.055, 0.056, 0.057, 0.059, 0.06, 0.061, 
    0.062, 0.063, 0.064, 0.065, 0.067, 0.068, 0.069, 0.071, 0.072, 0.073, 
    0.074, 0.075, 0.075, 0.076, 0.075, 0.075, 0.074, 0.073, 0.071, 0.069, 
    0.067, 0.065, 0.063, 0.061, 0.059, 0.057, 0.055, 0.053, 0.051, 0.049, 
    0.047, 0.046, 0.044, 0.043, 0.042, 0.041, 0.04, 0.039, 0.038, 0.037, 
    0.037, 0.036, 0.036, 0.036, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 
    0.035, 0.036, 0.036, 0.036, 0.036, 0.037, 0.037, 0.038, 0.038, 0.038, 
    0.038, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.038, 0.038, 0.037, 0.037, 0.036, 0.036, 0.035, 0.034, 
    0.034, 0.033, 0.032, 0.032, 0.031, 0.03, 0.029, 0.029, 0.028, 0.027, 
    0.026, 0.026, 0.025, 0.025, 0.024, 0.024, 0.023, 0.023, 0.022, 0.022, 
    0.021, 0.021, 0.02, 0.02, 0.02, 0.019, 0.019, 0.019, 0.018, 0.018, 0.018, 
    0.017, 0.017, 0.017, 0.016, 0.016, 0.016, 0.016, 0.015, 0.015, 0.015, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.013, 0.013, 0.013, 0.013, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.011, 0.011, 0.011, 0.011, 0.011, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.009, 0.009, 0.009, 0.009, 0.008, 0.008, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.013, 0.013, 0.013, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.014, 0.014, 0.014, 0.013, 0.013, 0.013, 0.013, 0.013, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.015, 0.015, 0.015, 0.015, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.017, 0.017, 0.017, 0.017, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.017, 0.017, 0.017, 0.017, 0.018, 0.018, 
    0.018, 0.019, 0.019, 0.02, 0.02, 0.021, 0.021, 0.022, 0.023, 0.023, 
    0.024, 0.025, 0.026, 0.026, 0.027, 0.028, 0.029, 0.03, 0.031, 0.032, 
    0.033, 0.034, 0.035, 0.037, 0.038, 0.039, 0.04, 0.041, 0.042, 0.043, 
    0.044, 0.044, 0.045, 0.046, 0.047, 0.048, 0.049, 0.05, 0.05, 0.051, 
    0.052, 0.053, 0.053, 0.054, 0.054, 0.055, 0.055, 0.056, 0.056, 0.057, 
    0.057, 0.057, 0.057, 0.058, 0.058, 0.058, 0.058, 0.058, 0.058, 0.059, 
    0.059, 0.059, 0.059, 0.059, 0.059, 0.059, 0.058, 0.058, 0.058, 0.058, 
    0.058, 0.057, 0.057, 0.057, 0.056, 0.055, 0.055, 0.054, 0.053, 0.052, 
    0.051, 0.05, 0.048, 0.047, 0.046, 0.045, 0.044, 0.042, 0.041, 0.04, 
    0.039, 0.038, 0.037, 0.036, 0.035, 0.034, 0.034, 0.033, 0.032, 0.032, 
    0.031, 0.03, 0.03, 0.029, 0.029, 0.029, 0.028, 0.028, 0.027, 0.027, 
    0.027, 0.026, 0.026, 0.026, 0.025, 0.025, 0.025, 0.024, 0.024, 0.024, 
    0.024, 0.023, 0.023, 0.023, 0.023, 0.022, 0.022, 0.022, 0.022, 0.021, 
    0.021, 0.021, 0.02, 0.02, 0.02, 0.02, 0.019, 0.019, 0.019, 0.018, 0.018, 
    0.018, 0.017, 0.017, 0.017, 0.017, 0.016, 0.016, 0.016, 0.016, 0.015, 
    0.015, 0.015, 0.015, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.009, 0.009, 0.009, 0.008, 0.008, 0.007, 0.007, 0.006, 0.005, 0.004, 
    0.004, 0.003, 0.002, 0.003, 0.004, 0.005, 0.006, 0.006, 0.007, 0.008, 
    0.008, 0.008, 0.009, 0.009, 0.009, 0.01, 0.01, 0.011, 0.011, 0.012, 
    0.013, 0.014, 0.015, 0.015, 0.016, 0.016, 0.017, 0.017, 0.017, 0.017, 
    0.017, 0.017, 0.017, 0.017, 0.018, 0.018, 0.017, 0.017, 0.017, 0.017, 
    0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.016, 0.017, 
    0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.016, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 
    0.015, 0.015, 0.015, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009 ;

 idx_rfr_illite_img_ee = 0.042, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 
    0.043, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.045, 0.045, 0.045, 
    0.046, 0.046, 0.046, 0.047, 0.047, 0.048, 0.048, 0.048, 0.049, 0.049, 
    0.05, 0.05, 0.051, 0.051, 0.051, 0.052, 0.052, 0.051, 0.051, 0.051, 
    0.051, 0.05, 0.05, 0.049, 0.049, 0.048, 0.048, 0.047, 0.046, 0.046, 
    0.045, 0.044, 0.044, 0.043, 0.042, 0.042, 0.041, 0.04, 0.04, 0.039, 
    0.038, 0.037, 0.037, 0.036, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 
    0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 
    0.035, 0.035, 0.035, 0.035, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 
    0.034, 0.033, 0.033, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 
    0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 
    0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.034, 0.035, 0.035, 
    0.035, 0.035, 0.035, 0.035, 0.035, 0.036, 0.036, 0.036, 0.036, 0.036, 
    0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 
    0.036, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 
    0.034, 0.034, 0.034, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 0.035, 
    0.035, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 
    0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.037, 0.038, 0.038, 
    0.038, 0.038, 0.038, 0.038, 0.038, 0.039, 0.039, 0.039, 0.039, 0.039, 
    0.039, 0.039, 0.04, 0.04, 0.04, 0.04, 0.04, 0.041, 0.041, 0.041, 0.041, 
    0.041, 0.041, 0.041, 0.041, 0.04, 0.04, 0.04, 0.04, 0.039, 0.039, 0.039, 
    0.039, 0.038, 0.038, 0.038, 0.037, 0.037, 0.037, 0.036, 0.036, 0.036, 
    0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.036, 0.037, 0.037, 
    0.037, 0.037, 0.037, 0.038, 0.038, 0.038, 0.038, 0.038, 0.038, 0.039, 
    0.039, 0.039, 0.039, 0.039, 0.039, 0.039, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.041, 0.041, 0.041, 0.041, 0.041, 0.042, 0.042, 0.042, 0.042, 0.042, 
    0.042, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.043, 0.044, 
    0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.045, 0.045, 0.045, 
    0.045, 0.045, 0.045, 0.046, 0.046, 0.046, 0.046, 0.047, 0.047, 0.047, 
    0.047, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 0.048, 
    0.048, 0.048, 0.048, 0.047, 0.047, 0.047, 0.047, 0.047, 0.046, 0.046, 
    0.046, 0.046, 0.046, 0.046, 0.045, 0.045, 0.045, 0.044, 0.044, 0.043, 
    0.043, 0.042, 0.042, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 0.041, 
    0.042, 0.042, 0.043, 0.044, 0.044, 0.045, 0.046, 0.047, 0.047, 0.048, 
    0.048, 0.048, 0.048, 0.048, 0.047, 0.047, 0.046, 0.046, 0.046, 0.045, 
    0.045, 0.045, 0.046, 0.046, 0.047, 0.048, 0.048, 0.049, 0.05, 0.051, 
    0.052, 0.052, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.053, 0.052, 
    0.052, 0.051, 0.051, 0.05, 0.05, 0.049, 0.048, 0.047, 0.047, 0.046, 
    0.046, 0.045, 0.045, 0.044, 0.044, 0.044, 0.044, 0.044, 0.044, 0.045, 
    0.045, 0.045, 0.046, 0.046, 0.046, 0.047, 0.047, 0.047, 0.047, 0.047, 
    0.047, 0.046, 0.046, 0.045, 0.045, 0.044, 0.044, 0.043, 0.042, 0.041, 
    0.04, 0.039, 0.037, 0.036, 0.034, 0.031, 0.029, 0.026, 0.023, 0.02, 
    0.017, 0.014, 0.011, 0.008, 0.005, 0.007, 0.009, 0.01, 0.011, 0.012, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.012, 0.012, 0.011, 0.011, 
    0.01, 0.01, 0.009, 0.008, 0.008, 0.007, 0.007, 0.006, 0.006, 0.005, 
    0.005, 0.004, 0.005, 0.005, 0.006, 0.006, 0.006, 0.007, 0.007, 0.007, 
    0.007, 0.007, 0.007, 0.006, 0.006, 0.006, 0.005, 0.005, 0.005, 0.005, 
    0.006, 0.006, 0.007, 0.008, 0.008, 0.009, 0.01, 0.01, 0.011, 0.011, 
    0.012, 0.012, 0.013, 0.013, 0.014, 0.014, 0.014, 0.014, 0.015, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.014, 0.013, 0.013, 0.013, 0.013, 0.013, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.007, 0.007, 
    0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 
    0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.008, 0.008, 0.008, 
    0.008, 0.009, 0.009, 0.009, 0.009, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.014, 0.014, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.015, 0.015, 0.015, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 
    0.015, 0.015, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.017, 0.017, 0.017, 
    0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 
    0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.016, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.017, 
    0.017, 0.017, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.015, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 
    0.015, 0.015, 0.016, 0.016, 0.016, 0.016, 0.016, 0.017, 0.017, 0.017, 
    0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.018, 0.018, 0.018, 0.018, 
    0.018, 0.018, 0.018, 0.018, 0.018, 0.018, 0.018, 0.018, 0.018, 0.018, 
    0.018, 0.018, 0.019, 0.019, 0.019, 0.019, 0.019, 0.019, 0.019, 0.019, 
    0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.021, 0.021, 0.021, 
    0.021, 0.021, 0.021, 0.021, 0.021, 0.022, 0.022, 0.022, 0.022, 0.022, 
    0.022, 0.022, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.026, 0.026, 0.026, 0.026, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 
    0.027, 0.028, 0.028, 0.028, 0.028, 0.028, 0.027, 0.027, 0.027, 0.027, 
    0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 
    0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.027, 0.028, 0.028, 0.028, 
    0.028, 0.028, 0.028, 0.029, 0.029, 0.029, 0.03, 0.03, 0.03, 0.03, 0.031, 
    0.031, 0.032, 0.032, 0.032, 0.033, 0.033, 0.034, 0.034, 0.035, 0.035, 
    0.036, 0.036, 0.037, 0.038, 0.038, 0.039, 0.039, 0.04, 0.04, 0.041, 
    0.042, 0.042, 0.043, 0.043, 0.044, 0.044, 0.045, 0.045, 0.045, 0.046, 
    0.046, 0.046, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.047, 0.046, 
    0.046, 0.046, 0.045, 0.045, 0.045, 0.044, 0.044, 0.043, 0.042, 0.042, 
    0.041, 0.04, 0.04, 0.039, 0.038, 0.037, 0.036, 0.035, 0.034, 0.033, 
    0.032, 0.031, 0.03, 0.029, 0.028, 0.027, 0.026, 0.024, 0.023, 0.022, 
    0.021, 0.02, 0.019, 0.018, 0.016, 0.015, 0.014, 0.013, 0.011, 0.01, 
    0.009, 0.007, 0.006, 0.005, 0.007, 0.008, 0.009, 0.011, 0.012, 0.013, 
    0.014, 0.015, 0.016, 0.017, 0.018, 0.019, 0.019, 0.02, 0.02, 0.02, 0.021, 
    0.021, 0.021, 0.021, 0.021, 0.021, 0.021, 0.02, 0.02, 0.02, 0.02, 0.02, 
    0.019, 0.019, 0.019, 0.019, 0.018, 0.018, 0.018, 0.018, 0.018, 0.018, 
    0.018, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 
    0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 0.016, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 
    0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.013, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.012, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.011, 0.011, 0.011, 0.012, 0.012, 0.012, 0.013, 0.013, 0.014, 0.015, 
    0.015, 0.016, 0.017, 0.017, 0.018, 0.018, 0.019, 0.02, 0.02, 0.021, 
    0.021, 0.022, 0.022, 0.023, 0.023, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 0.023, 
    0.023, 0.023, 0.023, 0.023, 0.023, 0.022, 0.022, 0.022, 0.021, 0.02, 
    0.02, 0.019, 0.019, 0.018, 0.018, 0.017, 0.017, 0.016, 0.016, 0.016, 
    0.015, 0.015, 0.015, 0.014, 0.014, 0.014, 0.014, 0.014, 0.014, 0.013, 
    0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.013, 0.012, 0.012, 0.012, 
    0.012, 0.012, 0.012, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.01, 0.009, 0.01, 0.009, 0.01, 
    0.009, 0.01, 0.009, 0.01, 0.009, 0.01, 0.009, 0.01, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.01, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.01, 0.01, 0.009, 0.01, 0.01, 0.009, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.011, 0.011, 0.011, 0.01, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 
    0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.011, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.008, 0.007, 0.006, 
    0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.005, 0.005, 0.004, 0.003, 
    0.002, 0.001, 0, 0, 0.001, 0.002, 0.002, 0.003, 0.003, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.003, 0.003, 0.003, 0.004, 0.004, 
    0.004, 0.005, 0.005, 0.005, 0.005, 0.006, 0.006, 0.006, 0.006, 0.006, 
    0.006, 0.006, 0.005, 0.005, 0.005, 0.005, 0.005, 0.004, 0.004, 0.004, 
    0.003, 0.003, 0.003, 0.002, 0.002, 0.002, 0.002, 0.003, 0.003, 0.003, 
    0.004, 0.005, 0.005, 0.005, 0.006, 0.007, 0.007, 0.007, 0.007, 0.007, 
    0.007, 0.006, 0.006, 0.006, 0.005, 0.004, 0.003, 0.002, 0.001, 0, 0.001, 
    0.001, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.002, 0.002, 0.002, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.003, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.005, 0.005, 0.005, 0.005, 0.005, 0.004, 0.004, 
    0.003, 0.003, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.003, 0.003, 
    0.004, 0.005, 0.005, 0.006, 0.006, 0.006, 0.007, 0.006, 0.005, 0.005, 
    0.004, 0.003, 0.003, 0.002, 0.002, 0.003, 0.004, 0.005, 0.006, 0.007, 
    0.009, 0.01, 0.01, 0.01, 0.01, 0.009, 0.008, 0.007, 0.006, 0.004, 0.003, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.003, 0.004, 0.004, 0.005, 
    0.005, 0.005, 0.005, 0.005, 0.004, 0.004, 0.004, 0.004, 0.005, 0.005, 
    0.006, 0.006, 0.007, 0.007, 0.007, 0.007, 0.007, 0.006, 0.006, 0.006, 
    0.005, 0.004, 0.004, 0.004, 0.004, 0.005, 0.005, 0.006, 0.006, 0.007, 
    0.008, 0.008, 0.008, 0.008, 0.008, 0.008, 0.007, 0.007, 0.006, 0.006, 
    0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 
    0.005, 0.005, 0.004, 0.004, 0.003, 0.003, 0.003, 0.003, 0.004, 0.004, 
    0.005, 0.005, 0.006, 0.007, 0.007, 0.008, 0.008, 0.007, 0.007, 0.007, 
    0.006, 0.006, 0.005, 0.005, 0.004, 0.004, 0.004, 0.004, 0.003, 0.003, 
    0.003, 0.003, 0.003, 0.004, 0.004, 0.004, 0.005, 0.005, 0.005, 0.006, 
    0.006, 0.006, 0.006, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 0.007, 
    0.007, 0.007, 0.008, 0.008, 0.008, 0.008, 0.008, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.01, 0.01, 0.01, 0.01, 0.01, 0.009, 0.009, 0.008, 0.008, 
    0.008, 0.007, 0.007, 0.007, 0.006, 0.006, 0.006, 0.005, 0.005, 0.005, 
    0.005, 0.005, 0.005, 0.005, 0.006, 0.006, 0.006, 0.006, 0.006, 0.006, 
    0.006, 0.006, 0.006, 0.006, 0.005, 0.005, 0.005, 0.004, 0.005, 0.004, 
    0.004, 0.004, 0.004 ;

 idx_rfr_illite_nr = 0.141, 0.141, 0.141, 0.142, 0.142, 0.142, 0.143, 0.143, 
    0.144, 0.145, 0.145, 0.146, 0.146, 0.147, 0.147, 0.148, 0.149, 0.15, 
    0.151, 0.152, 0.154, 0.155, 0.156, 0.157, 0.158, 0.16, 0.161, 0.162, 
    0.164, 0.165, 0.167, 0.167, 0.168, 0.169, 0.169, 0.169, 0.169, 0.168, 
    0.168, 0.168, 0.167, 0.166, 0.165, 0.164, 0.163, 0.162, 0.16, 0.159, 
    0.157, 0.156, 0.154, 0.153, 0.151, 0.149, 0.147, 0.145, 0.143, 0.14, 
    0.138, 0.135, 0.132, 0.129, 0.127, 0.125, 0.123, 0.123, 0.122, 0.122, 
    0.122, 0.122, 0.122, 0.121, 0.121, 0.121, 0.121, 0.121, 0.121, 0.12, 
    0.12, 0.12, 0.119, 0.119, 0.118, 0.117, 0.116, 0.116, 0.115, 0.115, 
    0.114, 0.114, 0.114, 0.114, 0.114, 0.114, 0.114, 0.114, 0.114, 0.114, 
    0.114, 0.115, 0.115, 0.115, 0.115, 0.115, 0.116, 0.116, 0.116, 0.116, 
    0.116, 0.116, 0.116, 0.115, 0.115, 0.115, 0.116, 0.116, 0.116, 0.117, 
    0.117, 0.118, 0.118, 0.119, 0.119, 0.12, 0.12, 0.121, 0.121, 0.122, 
    0.122, 0.122, 0.123, 0.123, 0.123, 0.122, 0.122, 0.121, 0.121, 0.12, 
    0.119, 0.119, 0.118, 0.118, 0.117, 0.117, 0.117, 0.116, 0.116, 0.116, 
    0.116, 0.116, 0.116, 0.116, 0.116, 0.117, 0.117, 0.117, 0.118, 0.119, 
    0.119, 0.12, 0.12, 0.121, 0.121, 0.121, 0.121, 0.122, 0.122, 0.122, 
    0.123, 0.123, 0.123, 0.124, 0.124, 0.125, 0.125, 0.126, 0.126, 0.126, 
    0.127, 0.127, 0.128, 0.128, 0.129, 0.129, 0.13, 0.13, 0.131, 0.132, 
    0.132, 0.133, 0.134, 0.134, 0.135, 0.136, 0.137, 0.137, 0.137, 0.138, 
    0.138, 0.138, 0.138, 0.138, 0.138, 0.137, 0.137, 0.137, 0.136, 0.135, 
    0.134, 0.133, 0.133, 0.132, 0.13, 0.129, 0.128, 0.127, 0.126, 0.125, 
    0.124, 0.123, 0.123, 0.123, 0.122, 0.122, 0.123, 0.123, 0.123, 0.124, 
    0.124, 0.125, 0.125, 0.126, 0.126, 0.127, 0.128, 0.128, 0.129, 0.129, 
    0.13, 0.13, 0.131, 0.131, 0.132, 0.132, 0.133, 0.133, 0.134, 0.134, 
    0.135, 0.136, 0.136, 0.137, 0.138, 0.138, 0.139, 0.14, 0.14, 0.141, 
    0.141, 0.142, 0.143, 0.143, 0.144, 0.144, 0.145, 0.145, 0.146, 0.146, 
    0.147, 0.147, 0.147, 0.148, 0.148, 0.149, 0.149, 0.15, 0.15, 0.151, 
    0.152, 0.152, 0.153, 0.153, 0.154, 0.155, 0.156, 0.156, 0.157, 0.158, 
    0.159, 0.16, 0.162, 0.163, 0.164, 0.165, 0.166, 0.167, 0.168, 0.168, 
    0.169, 0.169, 0.169, 0.169, 0.169, 0.169, 0.169, 0.169, 0.169, 0.169, 
    0.169, 0.169, 0.169, 0.169, 0.169, 0.169, 0.169, 0.169, 0.169, 0.168, 
    0.167, 0.166, 0.165, 0.163, 0.162, 0.16, 0.158, 0.156, 0.155, 0.154, 
    0.153, 0.153, 0.153, 0.154, 0.155, 0.156, 0.158, 0.161, 0.163, 0.166, 
    0.169, 0.171, 0.174, 0.175, 0.177, 0.177, 0.177, 0.177, 0.176, 0.175, 
    0.174, 0.172, 0.171, 0.171, 0.171, 0.171, 0.173, 0.174, 0.177, 0.179, 
    0.182, 0.185, 0.189, 0.192, 0.194, 0.197, 0.2, 0.202, 0.204, 0.206, 
    0.207, 0.208, 0.21, 0.211, 0.211, 0.212, 0.212, 0.213, 0.213, 0.212, 
    0.212, 0.212, 0.211, 0.21, 0.21, 0.209, 0.209, 0.208, 0.208, 0.208, 
    0.209, 0.209, 0.21, 0.212, 0.214, 0.216, 0.218, 0.221, 0.223, 0.226, 
    0.229, 0.232, 0.235, 0.238, 0.241, 0.244, 0.247, 0.25, 0.253, 0.256, 
    0.259, 0.263, 0.266, 0.27, 0.275, 0.279, 0.283, 0.288, 0.292, 0.297, 
    0.301, 0.304, 0.308, 0.31, 0.313, 0.314, 0.315, 0.315, 0.314, 0.312, 
    0.31, 0.307, 0.303, 0.298, 0.293, 0.287, 0.281, 0.274, 0.268, 0.261, 
    0.254, 0.247, 0.24, 0.234, 0.227, 0.221, 0.216, 0.211, 0.206, 0.202, 
    0.199, 0.195, 0.193, 0.19, 0.189, 0.187, 0.186, 0.186, 0.186, 0.187, 
    0.188, 0.189, 0.191, 0.193, 0.195, 0.197, 0.2, 0.203, 0.206, 0.208, 
    0.211, 0.214, 0.216, 0.219, 0.221, 0.223, 0.225, 0.228, 0.229, 0.231, 
    0.233, 0.234, 0.235, 0.236, 0.237, 0.238, 0.238, 0.238, 0.238, 0.237, 
    0.236, 0.235, 0.233, 0.231, 0.228, 0.226, 0.223, 0.22, 0.216, 0.213, 
    0.209, 0.206, 0.202, 0.198, 0.194, 0.19, 0.187, 0.183, 0.179, 0.176, 
    0.172, 0.168, 0.164, 0.161, 0.157, 0.153, 0.149, 0.145, 0.141, 0.138, 
    0.134, 0.13, 0.126, 0.122, 0.118, 0.114, 0.111, 0.107, 0.103, 0.0996, 
    0.0959, 0.0922, 0.0887, 0.0852, 0.0816, 0.0782, 0.0749, 0.0715, 0.0684, 
    0.0652, 0.0622, 0.0593, 0.0564, 0.0536, 0.051, 0.0485, 0.0461, 0.0439, 
    0.0417, 0.0397, 0.0378, 0.0361, 0.0345, 0.033, 0.0316, 0.0303, 0.0291, 
    0.0281, 0.0271, 0.0263, 0.0255, 0.0248, 0.0242, 0.0236, 0.0231, 0.0226, 
    0.0223, 0.022, 0.0217, 0.0215, 0.0214, 0.0214, 0.0214, 0.0214, 0.0214, 
    0.0215, 0.0215, 0.0216, 0.0216, 0.0216, 0.0216, 0.0216, 0.0215, 0.0214, 
    0.0214, 0.0213, 0.0212, 0.0212, 0.0211, 0.0211, 0.0211, 0.0211, 0.0212, 
    0.0212, 0.0213, 0.0214, 0.0214, 0.0215, 0.0216, 0.0217, 0.0218, 0.022, 
    0.0222, 0.0223, 0.0225, 0.0227, 0.0229, 0.0232, 0.0234, 0.0236, 0.0239, 
    0.0243, 0.0246, 0.0249, 0.0253, 0.0257, 0.026, 0.0265, 0.0268, 0.0271, 
    0.0276, 0.0279, 0.0282, 0.0286, 0.0289, 0.0291, 0.0294, 0.0297, 0.03, 
    0.0302, 0.0305, 0.0308, 0.031, 0.0313, 0.0316, 0.0319, 0.0322, 0.0325, 
    0.0327, 0.033, 0.0331, 0.0333, 0.0333, 0.0332, 0.0331, 0.0329, 0.0326, 
    0.0323, 0.032, 0.0316, 0.0314, 0.0312, 0.031, 0.0309, 0.0309, 0.031, 
    0.0312, 0.0314, 0.0317, 0.032, 0.0323, 0.0327, 0.0331, 0.0334, 0.0338, 
    0.0342, 0.0345, 0.0349, 0.0352, 0.0356, 0.036, 0.0364, 0.0367, 0.0371, 
    0.0375, 0.0378, 0.0382, 0.0384, 0.0388, 0.039, 0.0393, 0.0395, 0.0397, 
    0.04, 0.0402, 0.0406, 0.0409, 0.0413, 0.0416, 0.042, 0.0424, 0.0428, 
    0.0432, 0.0437, 0.0441, 0.0444, 0.0448, 0.0452, 0.0454, 0.0457, 0.0459, 
    0.046, 0.0461, 0.0461, 0.0461, 0.0461, 0.0461, 0.0461, 0.0461, 0.0461, 
    0.0461, 0.0462, 0.0463, 0.0464, 0.0465, 0.0468, 0.0471, 0.0474, 0.0479, 
    0.0483, 0.0488, 0.0494, 0.0498, 0.0503, 0.0507, 0.051, 0.0512, 0.0512, 
    0.0509, 0.0505, 0.05, 0.0494, 0.0486, 0.0478, 0.047, 0.0463, 0.0457, 
    0.0454, 0.0452, 0.0452, 0.0453, 0.0456, 0.046, 0.0464, 0.0468, 0.047, 
    0.047, 0.0468, 0.0465, 0.0458, 0.0449, 0.0439, 0.0426, 0.0413, 0.0402, 
    0.039, 0.038, 0.0372, 0.0367, 0.0364, 0.0365, 0.0368, 0.0373, 0.038, 
    0.0389, 0.0399, 0.0408, 0.0419, 0.0428, 0.0437, 0.0446, 0.0454, 0.0461, 
    0.0468, 0.0474, 0.0479, 0.0485, 0.0489, 0.0493, 0.0497, 0.05, 0.0503, 
    0.0505, 0.0508, 0.051, 0.0512, 0.0514, 0.0516, 0.0518, 0.052, 0.0523, 
    0.0525, 0.0529, 0.0532, 0.0536, 0.054, 0.0545, 0.055, 0.0555, 0.056, 
    0.0565, 0.0571, 0.0576, 0.0581, 0.0586, 0.0591, 0.0596, 0.06, 0.0606, 
    0.0611, 0.0616, 0.0621, 0.0627, 0.0632, 0.0637, 0.0642, 0.0648, 0.0653, 
    0.0658, 0.0664, 0.067, 0.0675, 0.068, 0.0685, 0.0691, 0.0697, 0.0702, 
    0.0708, 0.0714, 0.072, 0.0725, 0.0731, 0.0737, 0.0742, 0.0748, 0.0754, 
    0.0759, 0.0765, 0.0771, 0.0777, 0.0784, 0.079, 0.0798, 0.0806, 0.0813, 
    0.0822, 0.0832, 0.0842, 0.0851, 0.0861, 0.0871, 0.088, 0.0889, 0.0897, 
    0.0904, 0.0912, 0.0917, 0.0922, 0.0925, 0.0927, 0.0928, 0.0929, 0.0928, 
    0.0927, 0.0926, 0.0924, 0.0922, 0.0919, 0.0917, 0.0914, 0.0913, 0.0911, 
    0.091, 0.0909, 0.0909, 0.0909, 0.091, 0.0911, 0.0913, 0.0915, 0.0918, 
    0.0921, 0.0925, 0.0928, 0.0934, 0.0939, 0.0945, 0.0952, 0.0959, 0.0967, 
    0.0975, 0.0984, 0.0994, 0.101, 0.102, 0.103, 0.104, 0.105, 0.107, 0.108, 
    0.11, 0.111, 0.113, 0.115, 0.117, 0.119, 0.12, 0.122, 0.124, 0.127, 
    0.129, 0.131, 0.133, 0.135, 0.138, 0.14, 0.142, 0.145, 0.147, 0.149, 
    0.152, 0.154, 0.157, 0.159, 0.162, 0.164, 0.167, 0.17, 0.172, 0.175, 
    0.177, 0.179, 0.182, 0.184, 0.186, 0.189, 0.191, 0.193, 0.195, 0.197, 
    0.199, 0.201, 0.203, 0.205, 0.207, 0.209, 0.211, 0.213, 0.215, 0.217, 
    0.219, 0.221, 0.223, 0.225, 0.226, 0.228, 0.23, 0.232, 0.234, 0.235, 
    0.237, 0.239, 0.24, 0.242, 0.244, 0.246, 0.248, 0.25, 0.251, 0.254, 
    0.256, 0.258, 0.26, 0.262, 0.265, 0.268, 0.27, 0.273, 0.276, 0.279, 
    0.282, 0.285, 0.288, 0.29, 0.293, 0.296, 0.299, 0.301, 0.303, 0.305, 
    0.307, 0.308, 0.309, 0.31, 0.31, 0.31, 0.31, 0.309, 0.308, 0.307, 0.305, 
    0.303, 0.301, 0.299, 0.296, 0.293, 0.291, 0.288, 0.285, 0.282, 0.279, 
    0.276, 0.273, 0.27, 0.268, 0.265, 0.263, 0.26, 0.258, 0.256, 0.254, 
    0.252, 0.251, 0.249, 0.247, 0.245, 0.244, 0.242, 0.241, 0.239, 0.238, 
    0.237, 0.236, 0.235, 0.234, 0.233, 0.233, 0.232, 0.232, 0.231, 0.231, 
    0.231, 0.23, 0.23, 0.229, 0.229, 0.228, 0.227, 0.226, 0.225, 0.224, 
    0.222, 0.221, 0.219, 0.218, 0.216, 0.214, 0.212, 0.21, 0.208, 0.206, 
    0.204, 0.201, 0.199, 0.197, 0.195, 0.192, 0.19, 0.188, 0.186, 0.184, 
    0.181, 0.179, 0.177, 0.175, 0.173, 0.171, 0.168, 0.166, 0.164, 0.162, 
    0.16, 0.158, 0.156, 0.154, 0.151, 0.149, 0.147, 0.145, 0.142, 0.14, 
    0.137, 0.135, 0.132, 0.129, 0.127, 0.124, 0.121, 0.117, 0.114, 0.11, 
    0.106, 0.102, 0.0984, 0.0943, 0.0903, 0.0863, 0.0825, 0.079, 0.076, 
    0.0733, 0.0711, 0.0693, 0.0679, 0.0668, 0.0661, 0.0654, 0.0648, 0.0642, 
    0.0634, 0.0625, 0.0613, 0.06, 0.0584, 0.0567, 0.0547, 0.0527, 0.0507, 
    0.0485, 0.0465, 0.0445, 0.0426, 0.0408, 0.039, 0.0373, 0.0358, 0.0342, 
    0.0329, 0.0314, 0.0302, 0.0289, 0.0277, 0.0266, 0.0255, 0.0245, 0.0235, 
    0.0225, 0.0217, 0.0209, 0.0201, 0.0193, 0.0186, 0.0179, 0.0172, 0.0165, 
    0.0159, 0.0152, 0.0145, 0.0138, 0.0132, 0.0126, 0.0119, 0.0113, 0.0107, 
    0.0101, 0.0096, 0.0091, 0.0086, 0.00815, 0.00775, 0.00735, 0.00695, 
    0.00655, 0.00615, 0.0058, 0.00545, 0.0051, 0.0048, 0.00445, 0.0042, 
    0.0039, 0.00365, 0.0034, 0.0032, 0.003, 0.00285, 0.0027, 0.0026, 0.0025, 
    0.0024, 0.0023, 0.0022, 0.0021, 0.00205, 0.00195, 0.0019, 0.00185, 
    0.0018, 0.00175, 0.00175, 0.00175, 0.00175, 0.0018, 0.0018, 0.00185, 
    0.0019, 0.00195, 0.00195, 0.002, 0.00195, 0.00195, 0.00195, 0.0019, 
    0.0019, 0.00185, 0.0018, 0.0018, 0.0018, 0.0018, 0.00185, 0.00185, 
    0.0019, 0.002, 0.00205, 0.00215, 0.0022, 0.0023, 0.00235, 0.0024, 0.0025, 
    0.00255, 0.00265, 0.00275, 0.0028, 0.0029, 0.003, 0.0031, 0.0032, 0.0033, 
    0.0034, 0.0035, 0.00355, 0.0036, 0.00365, 0.0037, 0.0037, 0.00375, 
    0.00375, 0.0038, 0.00385, 0.0039, 0.004, 0.0041, 0.0042, 0.0043, 0.0044, 
    0.00455, 0.00465, 0.0047, 0.0048, 0.0049, 0.00495, 0.005, 0.00505, 
    0.0051, 0.00515, 0.0052, 0.00525, 0.0053, 0.00535, 0.00545, 0.0055, 
    0.00555, 0.0056, 0.00565, 0.0057, 0.00575, 0.0058, 0.00585, 0.00595, 
    0.006, 0.0061, 0.0062, 0.0063, 0.0064, 0.00645, 0.00655, 0.0066, 0.0067, 
    0.00675, 0.0068, 0.00685, 0.0069, 0.00695, 0.007, 0.00705, 0.0071, 
    0.00715, 0.00725, 0.0073, 0.0074, 0.00745, 0.00755, 0.00765, 0.0077, 
    0.0078, 0.00785, 0.00795, 0.008, 0.0081, 0.00815, 0.00825, 0.0083, 
    0.00835, 0.00845, 0.0085, 0.0086, 0.00865, 0.00875, 0.0088, 0.00885, 
    0.00895, 0.009, 0.00905, 0.00915, 0.0092, 0.00925, 0.0093, 0.0094, 
    0.00945, 0.0095, 0.00955, 0.0096, 0.0097, 0.00975, 0.0098, 0.00985, 
    0.0099, 0.00995, 0.01, 0.01, 0.0101, 0.0102, 0.0102, 0.0103, 0.0103, 
    0.0104, 0.0104, 0.0104, 0.0104, 0.0105, 0.0105, 0.0105, 0.0106, 0.0106, 
    0.0107, 0.0108, 0.0108, 0.0109, 0.0109, 0.011, 0.011, 0.011, 0.011, 
    0.0111, 0.0111, 0.0111, 0.0112, 0.0113, 0.0113, 0.0113, 0.0114, 0.0114, 
    0.0114, 0.0114, 0.0115, 0.0115, 0.0115, 0.0115, 0.0116, 0.0116, 0.0116, 
    0.0117, 0.0117, 0.0117, 0.0117, 0.0118, 0.0118, 0.0119, 0.0119, 0.0119, 
    0.0119, 0.012, 0.012, 0.012, 0.012, 0.0121, 0.0121, 0.0121, 0.0121, 
    0.0121, 0.0121, 0.0122, 0.0122, 0.0122, 0.0122, 0.0123, 0.0123, 0.0124, 
    0.0124, 0.0124, 0.0124, 0.0124, 0.0124, 0.0125, 0.0125, 0.0125, 0.0125, 
    0.0125, 0.0125, 0.0125, 0.0126, 0.0126, 0.0126, 0.0126, 0.0126, 0.0126, 
    0.0126, 0.0127, 0.0127, 0.0127, 0.0127, 0.0127, 0.0128, 0.0128, 0.0128, 
    0.0128, 0.0129, 0.0129, 0.013, 0.013, 0.013, 0.013, 0.013, 0.0131, 
    0.0131, 0.0131, 0.0131, 0.0131, 0.0131, 0.0131, 0.0132, 0.0132, 0.0132, 
    0.0132, 0.0132, 0.0132, 0.0132, 0.0133, 0.0133, 0.0133, 0.0133, 0.0134, 
    0.0134, 0.0135, 0.0135, 0.0135, 0.0135, 0.0136, 0.0136, 0.0136, 0.0136, 
    0.0136, 0.0137, 0.0137, 0.0137, 0.0137, 0.0137, 0.0138, 0.0138, 0.0138, 
    0.0138, 0.0139, 0.0139, 0.0139, 0.0139, 0.014, 0.014, 0.0141, 0.0141, 
    0.0141, 0.0141, 0.0141, 0.0142, 0.0142, 0.0142, 0.0143, 0.0143, 0.0143, 
    0.0143, 0.0143, 0.0144, 0.0144, 0.0144, 0.0144, 0.0145, 0.0146, 0.0146, 
    0.0146, 0.0146, 0.0147, 0.0147, 0.0147, 0.0148, 0.0148, 0.0148, 0.0148, 
    0.0148, 0.0149, 0.0149, 0.0149, 0.015, 0.015, 0.015, 0.015, 0.0151, 
    0.0152, 0.0152, 0.0152, 0.0152, 0.0153, 0.0153, 0.0153, 0.0154, 0.0154, 
    0.0154, 0.0154, 0.0154, 0.0155, 0.0155, 0.0155, 0.0156, 0.0156, 0.0157, 
    0.0157, 0.0157, 0.0158, 0.0158, 0.0158, 0.0158, 0.0159, 0.0159, 0.0159, 
    0.0159, 0.0159, 0.0159, 0.016, 0.016, 0.016, 0.016, 0.0161, 0.0161, 
    0.0161, 0.0162, 0.0162, 0.0162, 0.0162, 0.0163, 0.0163, 0.0163, 0.0163, 
    0.0164, 0.0164, 0.0165, 0.0165, 0.0165, 0.0166, 0.0166, 0.0166, 0.0166, 
    0.0167, 0.0167, 0.0167, 0.0167, 0.0168, 0.0168, 0.0168, 0.0168, 0.0169, 
    0.0169, 0.0169, 0.0169, 0.0169, 0.017, 0.017, 0.017, 0.017, 0.017, 0.017, 
    0.0171, 0.0171, 0.0171, 0.0171, 0.0172, 0.0172, 0.0172, 0.0172, 0.0172, 
    0.0172, 0.0172, 0.0173, 0.0173, 0.0173, 0.0173, 0.0173, 0.0173, 0.0174, 
    0.0174, 0.0174, 0.0174, 0.0174, 0.0175, 0.0175, 0.0176, 0.0176, 0.0176, 
    0.0176, 0.0176, 0.0176, 0.0177, 0.0177, 0.0177, 0.0177, 0.0177, 0.0177, 
    0.0177, 0.0178, 0.0178, 0.0178, 0.0178, 0.0178, 0.0179, 0.0179, 0.0179, 
    0.0179, 0.0179, 0.018, 0.018, 0.018, 0.018, 0.018, 0.018, 0.0181, 0.0181, 
    0.0181, 0.0181, 0.0181, 0.0181, 0.0181, 0.0181, 0.0181, 0.0182, 0.0182, 
    0.0182, 0.0182, 0.0182, 0.0182, 0.0183, 0.0183, 0.0183, 0.0183, 0.0183, 
    0.0183, 0.0183, 0.0184, 0.0184, 0.0184, 0.0184, 0.0184, 0.0184, 0.0184, 
    0.0184, 0.0184, 0.0185, 0.0185, 0.0185, 0.0185, 0.0185, 0.0186, 0.0186, 
    0.0186, 0.0187, 0.0187, 0.0187, 0.0187, 0.0187, 0.0187, 0.0188, 0.0188, 
    0.0188, 0.0188, 0.0188, 0.0188, 0.0188, 0.0189, 0.0189, 0.0189, 0.0189, 
    0.0189, 0.0189, 0.0189, 0.0189, 0.0189, 0.019, 0.019, 0.019, 0.019, 
    0.019, 0.019, 0.0191, 0.0191, 0.0191, 0.0191, 0.0191, 0.0191, 0.0191, 
    0.0191, 0.0191, 0.0192, 0.0192, 0.0192, 0.0192, 0.0192, 0.0192, 0.0192, 
    0.0192, 0.0192, 0.0192, 0.0193, 0.0193, 0.0193, 0.0193, 0.0193, 0.0193, 
    0.0193, 0.0193, 0.0194, 0.0194, 0.0194, 0.0194, 0.0194, 0.0194, 0.0194, 
    0.0194, 0.0195, 0.0195, 0.0195, 0.0195, 0.0195, 0.0195, 0.0195, 0.0195, 
    0.0196, 0.0196, 0.0196, 0.0196, 0.0196, 0.0196, 0.0197, 0.0197, 0.0197, 
    0.0197, 0.0197, 0.0197, 0.0197, 0.0197, 0.0197, 0.0197, 0.0198, 0.0198, 
    0.0198, 0.0198, 0.0198, 0.0198, 0.0198, 0.0198, 0.0198, 0.0198, 0.0199, 
    0.0199, 0.0199, 0.0199, 0.0199, 0.0199, 0.0199, 0.02, 0.02, 0.02, 0.02, 
    0.02, 0.02, 0.02, 0.02, 0.0201, 0.0201, 0.0201, 0.0201, 0.0201, 0.0201, 
    0.0201, 0.0201, 0.0201, 0.0201, 0.0202, 0.0202, 0.0202, 0.0202, 0.0202, 
    0.0203, 0.0203, 0.0203, 0.0203, 0.0203, 0.0203, 0.0203, 0.0203, 0.0203, 
    0.0203, 0.0203, 0.0203, 0.0203, 0.0203, 0.0203, 0.0203, 0.0203, 0.0203, 
    0.0203, 0.0203, 0.0204, 0.0204, 0.0204, 0.0204, 0.0204, 0.0204, 0.0204, 
    0.0204, 0.0204, 0.0204, 0.0205, 0.0205, 0.0205, 0.0205, 0.0205, 0.0205, 
    0.0205, 0.0205, 0.0206, 0.0206, 0.0206, 0.0206, 0.0206, 0.0206, 0.0206, 
    0.0207, 0.0207, 0.0207, 0.0207, 0.0207, 0.0207, 0.0207, 0.0207, 0.0207, 
    0.0207, 0.0208, 0.0208, 0.0208, 0.0209, 0.0209, 0.0209, 0.0209, 0.0209, 
    0.0209, 0.0209, 0.021, 0.021, 0.021, 0.021, 0.021, 0.021, 0.021, 0.021, 
    0.0211, 0.0211, 0.0211, 0.0211, 0.0211, 0.0211, 0.0211, 0.0212, 0.0212, 
    0.0212, 0.0212, 0.0212, 0.0212, 0.0212, 0.0212, 0.0212, 0.0212, 0.0213, 
    0.0213, 0.0213, 0.0213, 0.0213, 0.0213, 0.0214, 0.0214, 0.0214, 0.0214, 
    0.0214, 0.0214, 0.0214, 0.0214, 0.0214, 0.0215, 0.0215, 0.0215, 0.0215, 
    0.0215, 0.0215, 0.0216, 0.0216, 0.0216, 0.0216, 0.0216, 0.0216, 0.0216, 
    0.0217, 0.0217, 0.0217, 0.0217, 0.0217, 0.0217, 0.0217, 0.0218, 0.0218, 
    0.0218, 0.0218, 0.0218, 0.0218, 0.0218, 0.0218, 0.0219, 0.0219, 0.0219, 
    0.022, 0.022, 0.022, 0.022, 0.022, 0.022, 0.022, 0.0221, 0.0221, 0.0221, 
    0.0221, 0.0221, 0.0222, 0.0222, 0.0222, 0.0222, 0.0222, 0.0222, 0.0222, 
    0.0223, 0.0223, 0.0223, 0.0223, 0.0223, 0.0223, 0.0223, 0.0223, 0.0224, 
    0.0224, 0.0224, 0.0224, 0.0224, 0.0224, 0.0225, 0.0225, 0.0225, 0.0225, 
    0.0225, 0.0225, 0.0225, 0.0225, 0.0225, 0.0225, 0.0226, 0.0226, 0.0226, 
    0.0226, 0.0226, 0.0226, 0.0227, 0.0227, 0.0227, 0.0227, 0.0227, 0.0228, 
    0.0228, 0.0228, 0.0228, 0.0228, 0.0228, 0.0229, 0.0229, 0.0229, 0.0229, 
    0.0229, 0.0229, 0.0229, 0.0229, 0.0229, 0.023, 0.023, 0.023, 0.0231, 
    0.0231, 0.0231, 0.0231, 0.0231, 0.0231, 0.0232, 0.0232, 0.0232, 0.0232, 
    0.0232, 0.0232, 0.0232, 0.0233, 0.0233, 0.0233, 0.0233, 0.0233, 0.0233, 
    0.0233, 0.0233, 0.0233, 0.0234, 0.0234, 0.0234, 0.0234, 0.0234, 0.0234, 
    0.0234, 0.0234, 0.0234, 0.0234, 0.0235, 0.0235, 0.0235, 0.0235, 0.0235, 
    0.0235, 0.0235, 0.0235, 0.0235, 0.0235, 0.0236, 0.0236, 0.0236, 0.0236, 
    0.0236, 0.0236, 0.0236, 0.0236, 0.0236, 0.0236, 0.0236, 0.0236, 0.0236, 
    0.0236, 0.0236, 0.0237, 0.0237, 0.0237, 0.0237, 0.0237, 0.0237, 0.0237, 
    0.0237, 0.0237, 0.0237, 0.0238, 0.0238, 0.0238, 0.0238, 0.0238, 0.0238, 
    0.0238, 0.0238, 0.0238, 0.0238, 0.0239, 0.0239, 0.0239, 0.0239, 0.0239, 
    0.0239, 0.0239, 0.0239, 0.0239, 0.0239, 0.0239, 0.0239, 0.0239, 0.0239, 
    0.0239, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 
    0.024, 0.024, 0.024, 0.024, 0.024, 0.024, 0.0241, 0.0241, 0.0241, 0.0241, 
    0.0241, 0.0242, 0.0242, 0.0242, 0.0242, 0.0242, 0.0242, 0.0242, 0.0242, 
    0.0242, 0.0242, 0.0242, 0.0242, 0.0242, 0.0242, 0.0242, 0.0242, 0.0242, 
    0.0242, 0.0242, 0.0242, 0.0243, 0.0243, 0.0243, 0.0243, 0.0243, 0.0243, 
    0.0243, 0.0243, 0.0243, 0.0243, 0.0243, 0.0243, 0.0243, 0.0243, 0.0243, 
    0.0244, 0.0244, 0.0244, 0.0244, 0.0244, 0.0244, 0.0244, 0.0244, 0.0244, 
    0.0244, 0.0244, 0.0244, 0.0244, 0.0244, 0.0244, 0.0244, 0.0244, 0.0244, 
    0.0244, 0.0244, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 
    0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0246, 
    0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 
    0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 
    0.0246, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 
    0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 
    0.0247, 0.0247, 0.0247, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 
    0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 
    0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 
    0.0248, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 
    0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 
    0.0249, 0.0249, 0.0249, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.0251, 0.0251, 
    0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 
    0.0251, 0.0251, 0.0251, 0.0251, 0.0252, 0.0252, 0.0252, 0.0252, 0.0252, 
    0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 
    0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0254, 0.0254, 0.0254, 
    0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 
    0.0254, 0.0254, 0.0254, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 
    0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 
    0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 
    0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 
    0.0255, 0.0255, 0.0255, 0.0255, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 
    0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 
    0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 
    0.0255, 0.0255, 0.0255, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 
    0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 
    0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0257, 0.0257, 0.0257, 0.0257, 
    0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 
    0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 
    0.0257, 0.0257, 0.0257, 0.0257, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0256, 0.0255, 0.0255, 0.0255, 0.0255, 
    0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 
    0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 
    0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0255, 0.0254, 
    0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 
    0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 
    0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 
    0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 
    0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0253, 
    0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 
    0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 
    0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 
    0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 
    0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 
    0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 
    0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 
    0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 
    0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 0.0253, 
    0.0253, 0.0253, 0.0253, 0.0252, 0.0252, 0.0252, 0.0252, 0.0251, 0.0251, 
    0.0251, 0.0251, 0.0251, 0.0251, 0.0252, 0.0252, 0.0252, 0.0252, 0.0252, 
    0.0252, 0.0252, 0.0252, 0.0252, 0.0252, 0.0252, 0.0252, 0.0252, 0.0252, 
    0.0252, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 
    0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 
    0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 
    0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 
    0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 
    0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 
    0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.0251, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 
    0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 
    0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 
    0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 
    0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 
    0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 
    0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 
    0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 
    0.0249, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 
    0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 
    0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 
    0.0248, 0.0248, 0.0248, 0.0248, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 
    0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 
    0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 
    0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 
    0.0247, 0.0247, 0.0247, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 
    0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 
    0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 
    0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0245, 0.0245, 0.0245, 
    0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 
    0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 
    0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 
    0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 
    0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 
    0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 
    0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 0.0245, 
    0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 
    0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 
    0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 
    0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 
    0.0246, 0.0246, 0.0246, 0.0246, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 
    0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 
    0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 
    0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 
    0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0248, 
    0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0249, 0.0249, 
    0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0249, 0.0248, 0.0248, 
    0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 0.0247, 
    0.0248, 0.0249, 0.0249, 0.025, 0.025, 0.0251, 0.0251, 0.025, 0.025, 
    0.025, 0.0249, 0.0249, 0.0248, 0.0248, 0.0247, 0.0247, 0.0247, 0.0247, 
    0.0247, 0.0248, 0.0248, 0.0249, 0.025, 0.025, 0.0251, 0.0252, 0.0253, 
    0.0253, 0.0253, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0254, 0.0253, 
    0.0253, 0.0253, 0.0252, 0.0251, 0.0251, 0.025, 0.025, 0.0249, 0.0249, 
    0.0249, 0.0249, 0.0249, 0.025, 0.025, 0.0251, 0.0251, 0.0252, 0.0253, 
    0.0253, 0.0254, 0.0254, 0.0255, 0.0255, 0.0255, 0.0256, 0.0256, 0.0257, 
    0.0257, 0.0258, 0.0258, 0.0258, 0.0259, 0.0259, 0.0259, 0.026, 0.026, 
    0.026, 0.0259, 0.0259, 0.0259, 0.0258, 0.0258, 0.0257, 0.0256, 0.0255, 
    0.0254, 0.0253, 0.0252, 0.0251, 0.025, 0.025, 0.0249, 0.0249, 0.0249, 
    0.0248, 0.0248, 0.0248, 0.0248, 0.0248, 0.0247, 0.0247, 0.0246, 0.0245, 
    0.0244, 0.0242, 0.024, 0.0239, 0.0237, 0.0236, 0.0235, 0.0234, 0.0233, 
    0.0233, 0.0232, 0.0232, 0.0232, 0.0231, 0.0231, 0.0229, 0.0228, 0.0227, 
    0.0225, 0.0224, 0.0223, 0.0221, 0.022, 0.0218, 0.0217, 0.0216, 0.0215, 
    0.0215, 0.0215, 0.0215, 0.0215, 0.0216, 0.0216, 0.0217, 0.0218, 0.0218, 
    0.0219, 0.022, 0.022, 0.0219, 0.0218, 0.0218, 0.0217, 0.0216, 0.0215, 
    0.0214, 0.0214, 0.0214, 0.0214, 0.0214, 0.0214, 0.0214, 0.0215, 0.0216, 
    0.0217, 0.0218, 0.022, 0.0221, 0.0221, 0.0222, 0.0222, 0.0222, 0.0222, 
    0.0222, 0.0222, 0.0222, 0.0222, 0.0222, 0.0223, 0.0224, 0.0225, 0.0225, 
    0.0226, 0.0228, 0.0229, 0.0229, 0.0231, 0.0231, 0.0232, 0.0232, 0.0232, 
    0.0232, 0.0233, 0.0233, 0.0233, 0.0234, 0.0234, 0.0235, 0.0235, 0.0236, 
    0.0236, 0.0237, 0.0237, 0.0238, 0.0239, 0.024, 0.0241, 0.0242, 0.0243, 
    0.0243, 0.0244, 0.0244, 0.0245, 0.0245, 0.0246, 0.0246, 0.0246, 0.0247, 
    0.0247, 0.0247, 0.0247, 0.0247, 0.0246, 0.0246, 0.0246, 0.0246, 0.0246, 
    0.0246, 0.0246, 0.0247, 0.0247, 0.0247, 0.0248, 0.0249, 0.025, 0.0251, 
    0.0253, 0.0254, 0.0255, 0.0256, 0.0257, 0.0258, 0.0258, 0.0259, 0.0259, 
    0.0259, 0.0259, 0.0259, 0.0258, 0.0258, 0.0258, 0.0257, 0.0257, 0.0257, 
    0.0256, 0.0256, 0.0256, 0.0256, 0.0257, 0.0257, 0.0257, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0258, 0.0258, 0.0257, 0.0257, 0.0257, 0.0257, 0.0257, 
    0.0257, 0.0258, 0.0258, 0.0259, 0.026, 0.026, 0.0261, 0.0261, 0.0262, 
    0.0262, 0.0261, 0.0261, 0.026, 0.026, 0.0259, 0.0258, 0.0258, 0.0258, 
    0.0258, 0.0258, 0.0259, 0.026, 0.0261, 0.0262, 0.0264, 0.0265, 0.0265, 
    0.0264, 0.0264, 0.0262, 0.0261, 0.0259, 0.0258, 0.0256, 0.0255, 0.0254, 
    0.0254, 0.0254, 0.0255, 0.0256, 0.0258, 0.0258, 0.0259, 0.026, 0.0261, 
    0.0262, 0.0262, 0.0262, 0.0261, 0.0261, 0.0261, 0.0261, 0.0261, 0.0261, 
    0.0261, 0.0262, 0.0262, 0.0263, 0.0264, 0.0264, 0.0264, 0.0263, 0.0262, 
    0.0262, 0.0261, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.0261, 0.0262, 
    0.0263, 0.0264, 0.0264, 0.0264, 0.0264, 0.0264, 0.0264, 0.0263, 0.0262, 
    0.0261, 0.0261, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.0261, 
    0.0261, 0.0261, 0.0261, 0.0261, 0.026, 0.026, 0.026, 0.0259, 0.0259, 
    0.026, 0.026, 0.0261, 0.0261, 0.0262, 0.0263, 0.0264, 0.0265, 0.0265, 
    0.0265, 0.0265, 0.0265, 0.0264, 0.0264, 0.0262, 0.0262, 0.0261, 0.0261, 
    0.026, 0.026, 0.026, 0.026, 0.0261, 0.0261, 0.0261, 0.0262, 0.0262, 
    0.0263, 0.0264, 0.0264, 0.0265, 0.0265, 0.0266, 0.0266, 0.0266, 0.0266, 
    0.0266, 0.0266, 0.0266, 0.0266, 0.0266, 0.0266, 0.0266, 0.0266, 0.0266, 
    0.0266, 0.0266, 0.0266, 0.0266, 0.0266, 0.0266, 0.0266, 0.0266, 0.0265, 
    0.0265, 0.0265, 0.0265, 0.0265, 0.0264, 0.0264, 0.0264, 0.0263, 0.0262, 
    0.0262, 0.0261, 0.026, 0.026, 0.026, 0.0259, 0.0259, 0.0259, 0.0259, 
    0.0259, 0.0259, 0.026, 0.026, 0.026, 0.026, 0.0261, 0.0261, 0.0261, 
    0.0262, 0.0262, 0.0262, 0.0262, 0.0262, 0.0261, 0.0261, 0.0261, 0.0261, 
    0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 0.026, 
    0.026, 0.026 ;
}
